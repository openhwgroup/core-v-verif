`define  FORMAL  1

// TODO:silabs-robin  Re-enable core asserts.
`define  COREV_ASSERT_OFF  1
