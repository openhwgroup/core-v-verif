//
// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2020 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//


`ifndef __UVMT_CV32E40S_TB_SV__
`define __UVMT_CV32E40S_TB_SV__

/**
 * Module encapsulating the CV32E40S DUT wrapper, and associated SV interfaces.
 * Also provide UVM environment entry and exit points.
 */
`default_nettype none
module uvmt_cv32e40s_tb;

   import uvm_pkg::*;
   import cv32e40s_pkg::*;
   import uvmt_cv32e40s_pkg::*;
   import uvme_cv32e40s_pkg::*;
   `ifndef FORMAL
   import rvviApiPkg::*;
   `endif

   // Capture regs for test status from Virtual Peripheral in dut_wrap.mem_i
   bit        tp;
   bit        tf;
   bit        evalid;
   bit [31:0] evalue;

   // Agent interfaces
   uvma_isacov_if               isacov_if();
   uvma_clknrst_if              clknrst_if(); // clock and resets from the clknrst agent
   uvma_clknrst_if              clknrst_if_iss();
   uvma_debug_if                debug_if();
   uvma_interrupt_if            interrupt_if();
   uvma_clic_if                 clic_if();
   uvma_obi_memory_if #(
     .ADDR_WIDTH  (ENV_PARAM_INSTR_ADDR_WIDTH),
     .DATA_WIDTH  (ENV_PARAM_INSTR_DATA_WIDTH),
     .ACHK_WIDTH  (ENV_PARAM_INSTR_ACHK_WIDTH),
     .RCHK_WIDTH  (ENV_PARAM_INSTR_RCHK_WIDTH)
   ) obi_instr_if_i (
     .clk     (clknrst_if.clk),
     .reset_n (clknrst_if.reset_n)
   );

   uvma_obi_memory_if #(
     .ADDR_WIDTH  (ENV_PARAM_DATA_ADDR_WIDTH),
     .DATA_WIDTH  (ENV_PARAM_DATA_DATA_WIDTH),
     .ACHK_WIDTH  (ENV_PARAM_DATA_ACHK_WIDTH),
     .RCHK_WIDTH  (ENV_PARAM_DATA_RCHK_WIDTH)
   ) obi_data_if_i(
     .clk(clknrst_if.clk),
     .reset_n(clknrst_if.reset_n)
   );
   uvma_fencei_if               fencei_if_i(
     .clk(clknrst_if.clk),
     .reset_n(clknrst_if.reset_n)
   );

   // DUT Wrapper Interfaces
   uvmt_cv32e40s_vp_status_if       vp_status_if(.tests_passed(),
                                                 .tests_failed(),
                                                 .exit_valid(),
                                                 .exit_value()); // Status information generated by the Virtual Peripherals in the DUT WRAPPER memory.
   uvme_cv32e40s_core_cntrl_if      core_cntrl_if();
   uvmt_cv32e40s_core_status_if     core_status_if(.core_busy(),
                                                   .sec_lvl());     // Core status outputs

   // RVVI SystemVerilog Interface
   `ifndef FORMAL
      rvviTrace #( .NHART(1), .RETIRE(1)) rvvi_if();
   `endif

  /**
   * DUT WRAPPER instance:
   * This is an update of the riscv_wrapper.sv from PULP-Platform RI5CY project with
   * a few mods to bring unused ports from the CORE to this level using SV interfaces.
   */
   uvmt_cv32e40s_dut_wrap  #(
                             .B_EXT                (uvmt_cv32e40s_pkg::CORE_PARAM_B_EXT),
                             .DBG_NUM_TRIGGERS     (uvmt_cv32e40s_pkg::CORE_PARAM_DBG_NUM_TRIGGERS),
                             .DM_REGION_END        (uvmt_cv32e40s_pkg::CORE_PARAM_DM_REGION_END),
                             .DM_REGION_START      (uvmt_cv32e40s_pkg::CORE_PARAM_DM_REGION_START),
                             .LFSR0_CFG            (uvmt_cv32e40s_pkg::CORE_PARAM_LFSR0_CFG),
                             .LFSR1_CFG            (uvmt_cv32e40s_pkg::CORE_PARAM_LFSR1_CFG),
                             .LFSR2_CFG            (uvmt_cv32e40s_pkg::CORE_PARAM_LFSR2_CFG),
                             .M_EXT                (uvmt_cv32e40s_pkg::CORE_PARAM_M_EXT),
                             .PMA_CFG              (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_CFG),
                             .PMA_NUM_REGIONS      (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_NUM_REGIONS),
                             .PMP_GRANULARITY      (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_GRANULARITY),
                             .PMP_MSECCFG_RV       (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_MSECCFG_RV),
                             .PMP_NUM_REGIONS      (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_NUM_REGIONS),
                             .PMP_PMPADDR_RV       (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_PMPADDR_RV),
                             .PMP_PMPNCFG_RV       (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_PMPNCFG_RV),
                             .RV32                 (uvmt_cv32e40s_pkg::CORE_PARAM_RV32),
                             .SMCLIC               (uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC),
                             .SMCLIC_ID_WIDTH      (uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC_ID_WIDTH),
                             .SMCLIC_INTTHRESHBITS (uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC_INTTHRESHBITS),
                             .INSTR_ADDR_WIDTH     (ENV_PARAM_INSTR_ADDR_WIDTH),
                             .INSTR_RDATA_WIDTH    (ENV_PARAM_INSTR_DATA_WIDTH),
                             .RAM_ADDR_WIDTH       (ENV_PARAM_RAM_ADDR_WIDTH)
                            )
                            dut_wrap (
                              .clknrst_if(clknrst_if),
                              .interrupt_if(interrupt_if),
                              .vp_status_if(vp_status_if),
                              .core_cntrl_if(core_cntrl_if),
                              .core_status_if(core_status_if),
                              .obi_instr_if_i(obi_instr_if_i),
                              .obi_data_if_i(obi_data_if_i),
                              .fencei_if_i(fencei_if_i),
                              .clic_if(clic_if),
                              .*);

  bind cv32e40s_wrapper
    uvma_rvfi_instr_if#(uvme_cv32e40s_pkg::ILEN,
                        uvme_cv32e40s_pkg::XLEN) rvfi_instr_if_0_i(.clk(clk_i),
                                                                   .reset_n(rst_ni),

                                                                   .rvfi_valid(rvfi_i.rvfi_valid[0]),
                                                                   .rvfi_order(rvfi_i.rvfi_order[uvma_rvfi_pkg::ORDER_WL*0+:uvma_rvfi_pkg::ORDER_WL]),
                                                                   .rvfi_insn(rvfi_i.rvfi_insn[uvme_cv32e40s_pkg::ILEN*0+:uvme_cv32e40s_pkg::ILEN]),
                                                                   .rvfi_trap(rvfi_i.rvfi_trap),
                                                                   .rvfi_halt(rvfi_i.rvfi_halt[0]),
                                                                   .rvfi_intr(rvfi_i.rvfi_intr),
                                                                   .rvfi_dbg(rvfi_i.rvfi_dbg),
                                                                   .rvfi_dbg_mode(rvfi_i.rvfi_dbg_mode),
                                                                   .rvfi_nmip(rvfi_i.rvfi_nmip),
                                                                   .rvfi_mode(rvfi_i.rvfi_mode[uvma_rvfi_pkg::MODE_WL*0+:uvma_rvfi_pkg::MODE_WL]),
                                                                   .rvfi_ixl(rvfi_i.rvfi_ixl[uvma_rvfi_pkg::IXL_WL*0+:uvma_rvfi_pkg::IXL_WL]),
                                                                   .rvfi_pc_rdata(rvfi_i.rvfi_pc_rdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_pc_wdata(rvfi_i.rvfi_pc_wdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rs1_addr(rvfi_i.rvfi_rs1_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
                                                                   .rvfi_rs1_rdata(rvfi_i.rvfi_rs1_rdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rs2_addr(rvfi_i.rvfi_rs2_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
                                                                   .rvfi_rs2_rdata(rvfi_i.rvfi_rs2_rdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rs3_addr('0),
                                                                   .rvfi_rs3_rdata('0),
                                                                   .rvfi_rd1_addr(rvfi_i.rvfi_rd_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
                                                                   .rvfi_rd1_wdata(rvfi_i.rvfi_rd_wdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rd2_addr('0),
                                                                   .rvfi_rd2_wdata('0),
                                                                   .rvfi_gpr_rdata(rvfi_i.rvfi_gpr_rdata[32*uvme_cv32e40s_pkg::XLEN*0  +:32*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_gpr_rmask(rvfi_i.rvfi_gpr_rmask[32*0  +:32]),
                                                                   .rvfi_gpr_wdata(rvfi_i.rvfi_gpr_wdata[32*uvme_cv32e40s_pkg::XLEN*0  +:32*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_gpr_wmask(rvfi_i.rvfi_gpr_wmask[32*0  +:32]),
                                                                   .rvfi_mem_addr(rvfi_i.rvfi_mem_addr[  uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_mem_rdata(rvfi_i.rvfi_mem_rdata[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_mem_rmask(rvfi_i.rvfi_mem_rmask[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8*0  +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8]),
                                                                   .rvfi_mem_wdata(rvfi_i.rvfi_mem_wdata[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_mem_wmask(rvfi_i.rvfi_mem_wmask[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8*0  +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8])
                                                                   );

  // RVFI CSR binds
  `RVFI_CSR_BIND(cpuctrl)
  `RVFI_CSR_BIND(jvt)
  `RVFI_CSR_BIND(marchid)
  `RVFI_CSR_BIND(mcause)
  `RVFI_CSR_BIND(mcounteren)
  `RVFI_CSR_BIND(mcountinhibit)
  `RVFI_CSR_BIND(mcycle)
  `RVFI_CSR_BIND(mcycleh)
  `RVFI_CSR_BIND(menvcfg)
  `RVFI_CSR_BIND(menvcfgh)
  `RVFI_CSR_BIND(mepc)
  `RVFI_CSR_BIND(mhartid)
  `RVFI_CSR_BIND(mie)
  `RVFI_CSR_BIND(mimpid)
  `RVFI_CSR_BIND(minstret)
  `RVFI_CSR_BIND(minstreth)
  `RVFI_CSR_BIND(mip)
  `RVFI_CSR_BIND(misa)
  `RVFI_CSR_BIND(mscratch)
  `RVFI_CSR_BIND(mstateen0)
  `RVFI_CSR_BIND(mstateen1)
  `RVFI_CSR_BIND(mstateen2)
  `RVFI_CSR_BIND(mstateen3)
  `RVFI_CSR_BIND(mstateen0h)
  `RVFI_CSR_BIND(mstateen1h)
  `RVFI_CSR_BIND(mstateen2h)
  `RVFI_CSR_BIND(mstateen3h)
  `RVFI_CSR_BIND(mstatus)
  `RVFI_CSR_BIND(mstatush)
  `RVFI_CSR_BIND(mtval)
  `RVFI_CSR_BIND(mtvec)
  `RVFI_CSR_BIND(mvendorid)
  `RVFI_CSR_BIND(mseccfg)
  `RVFI_CSR_BIND(mseccfgh)

  `RVFI_CSR_BIND(dcsr)
  `RVFI_CSR_BIND(dpc)
  `RVFI_CSR_BIND(tselect)
  `RVFI_CSR_BIND(tinfo)
  `RVFI_CSR_BIND(tcontrol)

  `RVFI_CSR_IDX_BIND(mhpmcounter,,3)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,4)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,5)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,6)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,7)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,8)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,9)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,10)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,11)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,12)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,13)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,14)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,15)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,16)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,17)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,18)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,19)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,20)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,21)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,22)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,23)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,24)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,25)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,26)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,27)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,28)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,29)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,30)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,31)

  `RVFI_CSR_IDX_BIND(pmpcfg,,0)
  `RVFI_CSR_IDX_BIND(pmpcfg,,1)
  `RVFI_CSR_IDX_BIND(pmpcfg,,2)
  `RVFI_CSR_IDX_BIND(pmpcfg,,3)
  `RVFI_CSR_IDX_BIND(pmpcfg,,4)
  `RVFI_CSR_IDX_BIND(pmpcfg,,5)
  `RVFI_CSR_IDX_BIND(pmpcfg,,6)
  `RVFI_CSR_IDX_BIND(pmpcfg,,7)
  `RVFI_CSR_IDX_BIND(pmpcfg,,8)
  `RVFI_CSR_IDX_BIND(pmpcfg,,9)
  `RVFI_CSR_IDX_BIND(pmpcfg,,10)
  `RVFI_CSR_IDX_BIND(pmpcfg,,11)
  `RVFI_CSR_IDX_BIND(pmpcfg,,12)
  `RVFI_CSR_IDX_BIND(pmpcfg,,13)
  `RVFI_CSR_IDX_BIND(pmpcfg,,14)
  `RVFI_CSR_IDX_BIND(pmpcfg,,15)

  `RVFI_CSR_IDX_BIND(pmpaddr,,0)
  `RVFI_CSR_IDX_BIND(pmpaddr,,1)
  `RVFI_CSR_IDX_BIND(pmpaddr,,2)
  `RVFI_CSR_IDX_BIND(pmpaddr,,3)
  `RVFI_CSR_IDX_BIND(pmpaddr,,4)
  `RVFI_CSR_IDX_BIND(pmpaddr,,5)
  `RVFI_CSR_IDX_BIND(pmpaddr,,6)
  `RVFI_CSR_IDX_BIND(pmpaddr,,7)
  `RVFI_CSR_IDX_BIND(pmpaddr,,8)
  `RVFI_CSR_IDX_BIND(pmpaddr,,9)
  `RVFI_CSR_IDX_BIND(pmpaddr,,10)
  `RVFI_CSR_IDX_BIND(pmpaddr,,11)
  `RVFI_CSR_IDX_BIND(pmpaddr,,12)
  `RVFI_CSR_IDX_BIND(pmpaddr,,13)
  `RVFI_CSR_IDX_BIND(pmpaddr,,14)
  `RVFI_CSR_IDX_BIND(pmpaddr,,15)
  `RVFI_CSR_IDX_BIND(pmpaddr,,16)
  `RVFI_CSR_IDX_BIND(pmpaddr,,17)
  `RVFI_CSR_IDX_BIND(pmpaddr,,18)
  `RVFI_CSR_IDX_BIND(pmpaddr,,19)
  `RVFI_CSR_IDX_BIND(pmpaddr,,20)
  `RVFI_CSR_IDX_BIND(pmpaddr,,21)
  `RVFI_CSR_IDX_BIND(pmpaddr,,22)
  `RVFI_CSR_IDX_BIND(pmpaddr,,23)
  `RVFI_CSR_IDX_BIND(pmpaddr,,24)
  `RVFI_CSR_IDX_BIND(pmpaddr,,25)
  `RVFI_CSR_IDX_BIND(pmpaddr,,26)
  `RVFI_CSR_IDX_BIND(pmpaddr,,27)
  `RVFI_CSR_IDX_BIND(pmpaddr,,28)
  `RVFI_CSR_IDX_BIND(pmpaddr,,29)
  `RVFI_CSR_IDX_BIND(pmpaddr,,30)
  `RVFI_CSR_IDX_BIND(pmpaddr,,31)
  `RVFI_CSR_IDX_BIND(pmpaddr,,32)
  `RVFI_CSR_IDX_BIND(pmpaddr,,33)
  `RVFI_CSR_IDX_BIND(pmpaddr,,34)
  `RVFI_CSR_IDX_BIND(pmpaddr,,35)
  `RVFI_CSR_IDX_BIND(pmpaddr,,36)
  `RVFI_CSR_IDX_BIND(pmpaddr,,37)
  `RVFI_CSR_IDX_BIND(pmpaddr,,38)
  `RVFI_CSR_IDX_BIND(pmpaddr,,39)
  `RVFI_CSR_IDX_BIND(pmpaddr,,40)
  `RVFI_CSR_IDX_BIND(pmpaddr,,41)
  `RVFI_CSR_IDX_BIND(pmpaddr,,42)
  `RVFI_CSR_IDX_BIND(pmpaddr,,43)
  `RVFI_CSR_IDX_BIND(pmpaddr,,44)
  `RVFI_CSR_IDX_BIND(pmpaddr,,45)
  `RVFI_CSR_IDX_BIND(pmpaddr,,46)
  `RVFI_CSR_IDX_BIND(pmpaddr,,47)
  `RVFI_CSR_IDX_BIND(pmpaddr,,48)
  `RVFI_CSR_IDX_BIND(pmpaddr,,49)
  `RVFI_CSR_IDX_BIND(pmpaddr,,50)
  `RVFI_CSR_IDX_BIND(pmpaddr,,51)
  `RVFI_CSR_IDX_BIND(pmpaddr,,52)
  `RVFI_CSR_IDX_BIND(pmpaddr,,53)
  `RVFI_CSR_IDX_BIND(pmpaddr,,54)
  `RVFI_CSR_IDX_BIND(pmpaddr,,55)
  `RVFI_CSR_IDX_BIND(pmpaddr,,56)
  `RVFI_CSR_IDX_BIND(pmpaddr,,57)
  `RVFI_CSR_IDX_BIND(pmpaddr,,58)
  `RVFI_CSR_IDX_BIND(pmpaddr,,59)
  `RVFI_CSR_IDX_BIND(pmpaddr,,60)
  `RVFI_CSR_IDX_BIND(pmpaddr,,61)
  `RVFI_CSR_IDX_BIND(pmpaddr,,62)
  `RVFI_CSR_IDX_BIND(pmpaddr,,63)

  `RVFI_CSR_IDX_BIND(mhpmevent,,3)
  `RVFI_CSR_IDX_BIND(mhpmevent,,4)
  `RVFI_CSR_IDX_BIND(mhpmevent,,5)
  `RVFI_CSR_IDX_BIND(mhpmevent,,6)
  `RVFI_CSR_IDX_BIND(mhpmevent,,7)
  `RVFI_CSR_IDX_BIND(mhpmevent,,8)
  `RVFI_CSR_IDX_BIND(mhpmevent,,9)
  `RVFI_CSR_IDX_BIND(mhpmevent,,10)
  `RVFI_CSR_IDX_BIND(mhpmevent,,11)
  `RVFI_CSR_IDX_BIND(mhpmevent,,12)
  `RVFI_CSR_IDX_BIND(mhpmevent,,13)
  `RVFI_CSR_IDX_BIND(mhpmevent,,14)
  `RVFI_CSR_IDX_BIND(mhpmevent,,15)
  `RVFI_CSR_IDX_BIND(mhpmevent,,16)
  `RVFI_CSR_IDX_BIND(mhpmevent,,17)
  `RVFI_CSR_IDX_BIND(mhpmevent,,18)
  `RVFI_CSR_IDX_BIND(mhpmevent,,19)
  `RVFI_CSR_IDX_BIND(mhpmevent,,20)
  `RVFI_CSR_IDX_BIND(mhpmevent,,21)
  `RVFI_CSR_IDX_BIND(mhpmevent,,22)
  `RVFI_CSR_IDX_BIND(mhpmevent,,23)
  `RVFI_CSR_IDX_BIND(mhpmevent,,24)
  `RVFI_CSR_IDX_BIND(mhpmevent,,25)
  `RVFI_CSR_IDX_BIND(mhpmevent,,26)
  `RVFI_CSR_IDX_BIND(mhpmevent,,27)
  `RVFI_CSR_IDX_BIND(mhpmevent,,28)
  `RVFI_CSR_IDX_BIND(mhpmevent,,29)
  `RVFI_CSR_IDX_BIND(mhpmevent,,30)
  `RVFI_CSR_IDX_BIND(mhpmevent,,31)

  `RVFI_CSR_IDX_BIND(mhpmcounter,h,3)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,4)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,5)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,6)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,7)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,8)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,9)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,10)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,11)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,12)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,13)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,14)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,15)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,16)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,17)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,18)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,19)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,20)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,21)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,22)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,23)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,24)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,25)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,26)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,27)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,28)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,29)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,30)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,31)

  `RVFI_CSR_BIND(mconfigptr)
  `RVFI_CSR_BIND(secureseed0)
  `RVFI_CSR_BIND(secureseed1)
  `RVFI_CSR_BIND(secureseed2)

  if (CORE_PARAM_SMCLIC == 1) begin: gen_clic_rvfi_bind
    `RVFI_CSR_BIND(mintstatus)
    `RVFI_CSR_BIND(mintthresh)
    `RVFI_CSR_BIND(mnxti)
    `RVFI_CSR_BIND(mscratchcsw)
    `RVFI_CSR_BIND(mscratchcswl)
    `RVFI_CSR_BIND(mtvt)
  end : gen_clic_rvfi_bind

  // dscratch0
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_dscratch0_if_0_i(.clk(clk_i),
                                                                         .reset_n(rst_ni),
                                                                         .rvfi_csr_rmask(rvfi_i.rvfi_csr_dscratch_rmask[0]),
                                                                         .rvfi_csr_wmask(rvfi_i.rvfi_csr_dscratch_wmask[0]),
                                                                         .rvfi_csr_rdata(rvfi_i.rvfi_csr_dscratch_rdata[0]),
                                                                         .rvfi_csr_wdata(rvfi_i.rvfi_csr_dscratch_wdata[0])
    );

  // dscratch1
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_dscratch1_if_0_i(.clk(clk_i),
                                                                         .reset_n(rst_ni),
                                                                         .rvfi_csr_rmask(rvfi_i.rvfi_csr_dscratch_rmask[1]),
                                                                         .rvfi_csr_wmask(rvfi_i.rvfi_csr_dscratch_wmask[1]),
                                                                         .rvfi_csr_rdata(rvfi_i.rvfi_csr_dscratch_rdata[1]),
                                                                         .rvfi_csr_wdata(rvfi_i.rvfi_csr_dscratch_wdata[1])
    );

  // tdata1
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_tdata1_if_0_i(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[1]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[1]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[1]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[1])
    );

  // tdata2
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_tdata2_if_0_i(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[2]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[2]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[2]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[2])
    );

  // tdata3
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_tdata3_if_0_i(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[3]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[3]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[3]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[3])
    );

  bind cv32e40s_wrapper
    uvmt_cv32e40s_assumes  assumes_i (
      .obi  (dut_wrap.obi_instr_if_i),
      .rvfi (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i),
      .sup  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.support_logic_for_assert_coverage_modules_if),
      .*
    );

  bind uvmt_cv32e40s_dut_wrap
    uvma_obi_memory_assert_if_wrp#(
      .ADDR_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_ADDR_WIDTH),
      .DATA_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_DATA_WIDTH),
      .AUSER_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_AUSER_WIDTH),
      .WUSER_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_WUSER_WIDTH),
      .RUSER_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_RUSER_WIDTH),
      .ID_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_ID_WIDTH),
      .ACHK_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_ACHK_WIDTH),
      .RCHK_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_INSTR_RCHK_WIDTH),
      .IS_1P2(1)
    ) obi_instr_memory_assert_i(.obi(obi_instr_if_i));

  bind uvmt_cv32e40s_dut_wrap
    uvma_obi_memory_assert_if_wrp#(
      .ADDR_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_ADDR_WIDTH),
      .DATA_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_DATA_WIDTH),
      .AUSER_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_AUSER_WIDTH),
      .WUSER_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_WUSER_WIDTH),
      .RUSER_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_RUSER_WIDTH),
      .ID_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_ID_WIDTH),
      .ACHK_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_ACHK_WIDTH),
      .RCHK_WIDTH(uvme_cv32e40s_pkg::ENV_PARAM_DATA_RCHK_WIDTH),
      .IS_1P2(1)
    ) obi_data_memory_assert_i(.obi(obi_data_if_i));


  // Bind in verification modules to the design

  if (CORE_PARAM_SMCLIC == 0) begin: gen_interrupt_assert
    bind cv32e40s_core
      uvmt_cv32e40s_interrupt_assert  interrupt_assert_i (
        .mcause_n     ({cs_registers_i.mcause_n.irq, cs_registers_i.mcause_n.exception_code[4:0]}),
        .mip          (cs_registers_i.mip_rdata),
        .mie_q        (cs_registers_i.mie_q),
        .mstatus_mie  (cs_registers_i.mstatus_q.mie),
        .mstatus_tw   (cs_registers_i.mstatus_q.tw),
        .mtvec_mode_q (cs_registers_i.mtvec_q.mode),

        .if_stage_instr_req_o    (if_stage_i.m_c_obi_instr_if.s_req.req),
        .if_stage_instr_rvalid_i (if_stage_i.m_c_obi_instr_if.s_rvalid.rvalid),
        .if_stage_instr_rdata_i  (if_stage_i.m_c_obi_instr_if.resp_payload.rdata),
        .alignbuf_outstanding    (if_stage_i.prefetch_unit_i.alignment_buffer_i.outstanding_cnt_q),

        .ex_stage_instr_valid (ex_stage_i.id_ex_pipe_i.instr_valid),

        .wb_stage_instr_valid_i    (wb_stage_i.ex_wb_pipe_i.instr_valid),
        .wb_stage_instr_rdata_i    (wb_stage_i.ex_wb_pipe_i.instr.bus_resp.rdata),
        .wb_stage_instr_err_i      (wb_stage_i.ex_wb_pipe_i.instr.bus_resp.err),
        .wb_stage_instr_mpu_status (wb_stage_i.ex_wb_pipe_i.instr.mpu_status),

        .branch_taken_ex (controller_i.controller_fsm_i.branch_taken_ex),
        .debug_mode_q    (controller_i.controller_fsm_i.debug_mode_q),

        .irq_ack_o (core_i.irq_ack),
        .irq_id_o  (core_i.irq_id),

        .*
      );
  end : gen_interrupt_assert

  if (CORE_PARAM_SMCLIC == 1) begin: gen_clic_assert
    // CLIC assertions
    bind cv32e40s_core
      uvmt_cv32e40s_clic_interrupt_assert#(
        .SMCLIC (uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC)
      ) clic_assert_i(
        .dpc                 (cs_registers_i.dpc_rdata),
        .mintstatus          (cs_registers_i.mintstatus_rdata),
        .mintthresh          (cs_registers_i.mintthresh_rdata),
        .mcause              (cs_registers_i.mcause_rdata),
        .mtvec               (cs_registers_i.mtvec_rdata),
        .mtvt                (cs_registers_i.mtvt_rdata),
        .mepc                (cs_registers_i.mepc_rdata),
        .mip                 (cs_registers_i.mip_rdata),
        .mie                 (cs_registers_i.mie_rdata),
        .mnxti               (cs_registers_i.mnxti_rdata),
        .mscratch            (cs_registers_i.mscratch_rdata),
        .mscratchcsw         (cs_registers_i.mscratchcsw_rdata),
        .mscratchcswl        (cs_registers_i.mscratchcswl_rdata),
        .dcsr                (cs_registers_i.dcsr_rdata),

        .rvfi_mepc_wdata     (rvfi_i.rvfi_csr_mepc_wdata),
        .rvfi_mepc_wmask     (rvfi_i.rvfi_csr_mepc_wmask),
        .rvfi_mepc_rdata     (rvfi_i.rvfi_csr_mepc_rdata),
        .rvfi_mepc_rmask     (rvfi_i.rvfi_csr_mepc_rmask),
        .rvfi_dpc_rdata      (rvfi_i.rvfi_csr_dpc_rdata),
        .rvfi_dpc_rmask      (rvfi_i.rvfi_csr_dpc_rmask),
        .rvfi_mscratch_rdata (rvfi_i.rvfi_csr_mscratch_rdata),
        .rvfi_mscratch_rmask (rvfi_i.rvfi_csr_mscratch_rmask),
        .rvfi_mscratch_wdata (rvfi_i.rvfi_csr_mscratch_wdata),
        .rvfi_mscratch_wmask (rvfi_i.rvfi_csr_mscratch_wmask),
        .rvfi_mcause_wdata   (rvfi_i.rvfi_csr_mcause_wdata),
        .rvfi_mcause_wmask   (rvfi_i.rvfi_csr_mcause_wmask),

        .irq_i               (core_i.irq_i),
        .irq_ack             (core_i.irq_ack),
        .fetch_enable        (core_i.fetch_enable),
        .current_priv_mode   (core_i.priv_lvl),
        .mtvec_addr_i        (core_i.mtvec_addr_i),
        // External inputs
        .clic_if             (dut_wrap.clic_if),
        // Internal sampled   variants
        .irq_id              (core_i.irq_id[SMCLIC_ID_WIDTH-1:0]),
        .irq_level           (core_i.irq_level),
        .irq_priv            (core_i.irq_priv),
        .irq_shv             (core_i.irq_shv),

        .obi_instr_req       (core_i.instr_req_o),
        .obi_instr_gnt       (core_i.instr_gnt_i),
        .obi_instr_rvalid    (core_i.instr_rvalid_i),
        .obi_instr_addr      (core_i.instr_addr_o),
        .obi_instr_rdata     (core_i.instr_rdata_i),
        .obi_instr_rready    (1'b1),
        .obi_instr_err       (core_i.instr_err_i),

        .obi_data_addr       (core_i.data_addr_o),
        .obi_data_wdata      (core_i.data_wdata_o),
        .obi_data_we         (core_i.data_we_o),
        .obi_data_be         (core_i.data_be_o),
        .obi_data_req        (core_i.data_req_o),
        .obi_data_gnt        (core_i.data_gnt_i),
        .obi_data_rvalid     (core_i.data_rvalid_i),
        .obi_data_rready     (1'b1),
        .obi_data_err        (core_i.data_err_i),

        .debug_mode          (controller_i.controller_fsm_i.debug_mode_q),
        .debug_req           (core_i.debug_req_i),
        .debug_havereset     (core_i.debug_havereset_o),
        .debug_running       (core_i.debug_running_o),
        .debug_halt_addr     (dut_wrap.cv32e40s_wrapper_i.dm_halt_addr_i),
        .debug_exc_addr      (dut_wrap.cv32e40s_wrapper_i.dm_exception_addr_i),

        .rvfi_mode           (rvfi_i.rvfi_mode),
        .rvfi_insn           (rvfi_i.rvfi_insn),
        .rvfi_intr           (rvfi_i.rvfi_intr),
        .rvfi_rs1_rdata      (rvfi_i.rvfi_rs1_rdata),
        .rvfi_rs2_rdata      (rvfi_i.rvfi_rs2_rdata),
        .rvfi_rd_wdata       (rvfi_i.rvfi_rd_wdata),
        .rvfi_valid          (rvfi_i.rvfi_valid),
        .rvfi_pc_rdata       (rvfi_i.rvfi_pc_rdata),
        .rvfi_pc_wdata       (rvfi_i.rvfi_pc_wdata),
        .rvfi_trap           (rvfi_i.rvfi_trap),
        .rvfi_dbg_mode       (rvfi_i.rvfi_dbg_mode),
        .rvfi_dbg            (rvfi_i.rvfi_dbg),

        .wu_wfe              (dut_wrap.cv32e40s_wrapper_i.wu_wfe_i),
        .core_sleep_o        (core_i.core_sleep_o),
        .*
      );
  end : gen_clic_assert


  // User-mode assertions

  bind  cv32e40s_wrapper
    uvmt_cv32e40s_umode_assert  umode_assert_i (
      .rvfi_valid    (rvfi_i.rvfi_valid),
      .rvfi_mode     (rvfi_i.rvfi_mode),
      .rvfi_order    (rvfi_i.rvfi_order),
      .rvfi_trap     (rvfi_i.rvfi_trap),
      .rvfi_intr     (rvfi_i.rvfi_intr),
      .rvfi_insn     (rvfi_i.rvfi_insn),
      .rvfi_dbg_mode (rvfi_i.rvfi_dbg_mode),
      .rvfi_dbg      (rvfi_i.rvfi_dbg),
      .rvfi_pc_rdata (rvfi_i.rvfi_pc_rdata),

      .rvfi_csr_dcsr_rdata       (rvfi_i.rvfi_csr_dcsr_rdata),
      .rvfi_csr_mcause_rdata     (rvfi_i.rvfi_csr_mcause_rdata),
      .rvfi_csr_mcause_wdata     (rvfi_i.rvfi_csr_mcause_wdata),
      .rvfi_csr_mcause_wmask     (rvfi_i.rvfi_csr_mcause_wmask),
      .rvfi_csr_mcounteren_rdata (rvfi_i.rvfi_csr_mcounteren_rdata),
      .rvfi_csr_mie_rdata        (rvfi_i.rvfi_csr_mie_rdata),
      .rvfi_csr_mip_rdata        (rvfi_i.rvfi_csr_mip_rdata),
      .rvfi_csr_misa_rdata       (rvfi_i.rvfi_csr_misa_rdata),
      .rvfi_csr_mscratch_rdata   (rvfi_i.rvfi_csr_mscratch_rdata),
      .rvfi_csr_mscratch_rmask   (rvfi_i.rvfi_csr_mscratch_rmask),
      .rvfi_csr_mscratch_wdata   (rvfi_i.rvfi_csr_mscratch_wdata),
      .rvfi_csr_mscratch_wmask   (rvfi_i.rvfi_csr_mscratch_wmask),
      .rvfi_csr_mstateen0_rdata  (rvfi_i.rvfi_csr_mstateen0_rdata),
      .rvfi_csr_mstatus_rdata    (rvfi_i.rvfi_csr_mstatus_rdata),
      .rvfi_csr_mstatus_wdata    (rvfi_i.rvfi_csr_mstatus_wdata),
      .rvfi_csr_mstatus_wmask    (rvfi_i.rvfi_csr_mstatus_wmask),

      .mpu_iside_valid (core_i.if_stage_i.mpu_i.core_trans_valid_i),
      .mpu_iside_addr  (core_i.if_stage_i.mpu_i.core_trans_i.addr),

      .obi_iside_prot (core_i.instr_prot_o),
      .obi_dside_prot (core_i.data_prot_o),

      .*
    );


  // User-mode Coverage

  bind  cv32e40s_wrapper
    uvmt_cv32e40s_umode_cov  umode_cov_i (
      .rvfi_valid     (rvfi_i.rvfi_valid),
      .rvfi_trap      (rvfi_i.rvfi_trap),
      .rvfi_intr      (rvfi_i.rvfi_intr),
      .rvfi_insn      (rvfi_i.rvfi_insn),
      .rvfi_rs1_rdata (rvfi_i.rvfi_rs1_rdata),
      .rvfi_pc_rdata  (rvfi_i.rvfi_pc_rdata),
      .rvfi_mode      (rvfi_i.rvfi_mode),
      .rvfi_rd_addr   (rvfi_i.rvfi_rd_addr),
      .rvfi_dbg_mode  (rvfi_i.rvfi_dbg_mode),
      .rvfi_order     (rvfi_i.rvfi_order),
      .rvfi_mem_rmask (rvfi_i.rvfi_mem_rmask),
      .rvfi_mem_wmask (rvfi_i.rvfi_mem_wmask),

      .rvfi_csr_mstatus_rdata (rvfi_i.rvfi_csr_mstatus_rdata),
      .rvfi_csr_mstatus_rmask (rvfi_i.rvfi_csr_mstatus_rmask),
      .rvfi_csr_dcsr_rdata    (rvfi_i.rvfi_csr_dcsr_rdata),
      .rvfi_csr_dcsr_rmask    (rvfi_i.rvfi_csr_dcsr_rmask),

      .obi_iside_req  (core_i.instr_req_o),
      .obi_iside_gnt  (core_i.instr_gnt_i),
      .obi_iside_addr (core_i.instr_addr_o),
      .obi_iside_prot (core_i.instr_prot_o),

      .*
    );


  // Fence.i assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_fencei_assert #(
      .PMA_NUM_REGIONS (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_NUM_REGIONS),
      .PMA_CFG         (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_CFG)
    ) fencei_assert_i (
      .wb_valid           (core_i.wb_stage_i.wb_valid),
      .wb_instr_valid     (core_i.ex_wb_pipe.instr_valid),
      .wb_sys_en          (core_i.ex_wb_pipe.sys_en),
      .wb_sys_fencei_insn (core_i.ex_wb_pipe.sys_fencei_insn),
      .wb_pc              (core_i.ex_wb_pipe.pc),
      .wb_rdata           (core_i.ex_wb_pipe.instr.bus_resp.rdata),
      .wb_buffer_state    (core_i.load_store_unit_i.write_buffer_i.state),

      .rvfi_valid         (rvfi_i.rvfi_valid),
      .rvfi_intr          (rvfi_i.rvfi_intr.intr),
      .rvfi_dbg_mode      (rvfi_i.rvfi_dbg_mode),
      .rvfi_insn          (rvfi_i.rvfi_insn),

      .*
    );


  // RVFI assertions

  bind  dut_wrap.cv32e40s_wrapper_i.rvfi_i
    uvmt_cv32e40s_rvfi_assert #(
      .SMCLIC          (uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC),
      .SMCLIC_ID_WIDTH (uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC_ID_WIDTH)
    ) rvfi_assert_i (
      .rvfi             (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i),
      .writebuf_ready_o (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.ready_o),
      .writebuf_valid_i (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.valid_i),
      .*
    );


  // Core integration assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_integration_assert  integration_assert_i (.*);

  localparam PMP_ADDR_WIDTH = (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_GRANULARITY > 0) ? 33 - uvmt_cv32e40s_pkg::CORE_PARAM_PMP_GRANULARITY : 32;

  // Shadow:
  mseccfg_t pmp_mseccfg_q_shadow_q;
  pmpncfg_t pmpncfg_q_shadow_q[PMP_MAX_REGIONS];
  logic [PMP_ADDR_WIDTH-1:0] pmp_addr_q_shadow_q[PMP_MAX_REGIONS];

  mtvt_t mtvt_q_shadow_q;
  mtvec_t mtvec_q_shadow_q;
  mintstatus_t mintstatus_q_shadow_q;
  logic [31:0] mintthresh_q_shadow_q;
  logic [31:0] mie_q_hardened_shadow_q;

  // PMP register
  generate
    if (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_NUM_REGIONS > 0) begin
      assign pmp_mseccfg_q_shadow_q = (dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.csr_pmp.pmp_mseccfg_csr_i.gen_hardened.shadow_q);
    end else begin
      assign pmp_mseccfg_q_shadow_q = '0;
    end
  endgenerate

  generate for (genvar n = 0; n < uvmt_cv32e40s_pkg::CORE_PARAM_PMP_NUM_REGIONS; n++) begin
    assign pmpncfg_q_shadow_q[n] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.csr_pmp.gen_pmp_csr[n].pmp_region.pmpncfg_csr_i.gen_hardened.shadow_q;
    assign pmp_addr_q_shadow_q[n] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.csr_pmp.gen_pmp_csr[n].pmp_region.pmp_addr_csr_i.gen_hardened.shadow_q;
  end endgenerate

  generate
    if (SMCLIC==1) begin

      assign mtvt_q_shadow_q       = (dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.smclic_csrs.mtvt_csr_i.gen_hardened.shadow_q);
      assign mtvec_q_shadow_q      = (dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.smclic_csrs.mtvec_csr_i.gen_hardened.shadow_q);
      assign mintstatus_q_shadow_q = (dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.smclic_csrs.mintstatus_csr_i.gen_hardened.shadow_q);
      assign mintthresh_q_shadow_q = (dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.smclic_csrs.mintthresh_csr_i.gen_hardened.shadow_q);

      assign mie_q_hardened_shadow_q = '0;

    end else begin

      assign mtvt_q_shadow_q       = '0;
      assign mtvec_q_shadow_q      = (dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.basic_mode_csrs.mtvec_csr_i.gen_hardened.shadow_q);
      assign mintstatus_q_shadow_q = '0;
      assign mintthresh_q_shadow_q = '0;

      assign mie_q_hardened_shadow_q = (dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.basic_mode_csrs.mie_csr_i.gen_hardened.shadow_q);

    end
  endgenerate

  bind cv32e40s_wrapper
    uvmt_cv32e40s_xsecure_if
    #(.MTVT_ADDR_WIDTH   (core_i.MTVT_ADDR_WIDTH),
      .PMP_NUM_REGIONS   (PMP_NUM_REGIONS),
      .PMP_ADDR_WIDTH    (core_i.cs_registers_i.PMP_ADDR_WIDTH))

    xsecure_if (

      .core_i_sleep_unit_i_core_clock_gate_i_clk_en                                                                     (core_i.sleep_unit_i.core_clock_gate_i.clk_en),

      .core_i_data_err_i                                                                                                (core_i.data_err_i),
      .core_rf_we_wb                                                                                                    (core_i.rf_we_wb),
      .core_rf_waddr_wb                                                                                                 (core_i.rf_waddr_wb),
      .core_rf_wdata_wb                                                                                                 (core_i.rf_wdata_wb),
      .core_register_file_wrapper_register_file_mem                                                                     (core_i.register_file_wrapper_i.register_file_i.mem),
      .core_i_jump_target_id                                                                                            (core_i.jump_target_id),

      // OBI interface
      .core_i_if_stage_i_bus_resp                                                                                       (core_i.if_stage_i.bus_resp),
      .core_i_load_store_unit_i_bus_resp                                                                                (core_i.load_store_unit_i.bus_resp),

      .core_i_m_c_obi_data_if_req_payload                                                                               (core_i.m_c_obi_data_if.req_payload),
      .core_i_m_c_obi_data_if_resp_payload                                                                              (core_i.m_c_obi_data_if.resp_payload),
      .core_i_m_c_obi_instr_if_req_payload                                                                              (core_i.m_c_obi_instr_if.req_payload),
      .core_i_m_c_obi_instr_if_resp_payload                                                                             (core_i.m_c_obi_instr_if.resp_payload),

      .core_i_m_c_obi_data_if_s_req_req                                                                                 (core_i.m_c_obi_data_if.s_req.req),
      .core_i_m_c_obi_data_if_s_req_reqpar                                                                              (core_i.m_c_obi_data_if.s_req.reqpar),
      .core_i_m_c_obi_data_if_s_gnt_gnt                                                                                 (core_i.m_c_obi_data_if.s_gnt.gnt),
      .core_i_m_c_obi_data_if_s_gnt_gntpar                                                                              (core_i.m_c_obi_data_if.s_gnt.gntpar),
      .core_i_m_c_obi_data_if_s_rvalid_rvalid                                                                           (core_i.m_c_obi_data_if.s_rvalid.rvalid),
      .core_i_m_c_obi_data_if_s_rvalid_rvalidpar                                                                        (core_i.m_c_obi_data_if.s_rvalid.rvalidpar),

      .core_i_m_c_obi_instr_if_s_req_req                                                                                (core_i.m_c_obi_instr_if.s_req.req),
      .core_i_m_c_obi_instr_if_s_req_reqpar                                                                             (core_i.m_c_obi_instr_if.s_req.reqpar),
      .core_i_m_c_obi_instr_if_s_gnt_gnt                                                                                (core_i.m_c_obi_instr_if.s_gnt.gnt),
      .core_i_m_c_obi_instr_if_s_gnt_gntpar                                                                             (core_i.m_c_obi_instr_if.s_gnt.gntpar),
      .core_i_m_c_obi_instr_if_s_rvalid_rvalid                                                                          (core_i.m_c_obi_instr_if.s_rvalid.rvalid),
      .core_i_m_c_obi_instr_if_s_rvalid_rvalidpar                                                                       (core_i.m_c_obi_instr_if.s_rvalid.rvalidpar),

      .core_i_if_stage_i_prefetch_resp_valid                                                                            (core_i.if_stage_i.prefetch_resp_valid),
      .core_i_load_store_unit_i_resp_valid                                                                              (core_i.load_store_unit_i.resp_valid),
      .core_i_load_store_unit_i_bus_resp_valid                                                                          (core_i.load_store_unit_i.bus_resp_valid),

      .core_i_load_store_unit_i_response_filter_i_core_cnt_q                                                            (core_i.load_store_unit_i.response_filter_i.core_cnt_q),

      // CSR
      .core_alert_minor_o                                                                                               (core_i.alert_minor_o),
      .core_alert_major_o                                                                                               (core_i.alert_major_o),

      .core_xsecure_ctrl_cpuctrl_dataindtiming	                                                                        (core_i.xsecure_ctrl.cpuctrl.dataindtiming),
      .core_xsecure_ctrl_cpuctrl_rnddummy		                                                                            (core_i.xsecure_ctrl.cpuctrl.rnddummy),
      .core_xsecure_ctrl_cpuctrl_integrity                                                                              (core_i.xsecure_ctrl.cpuctrl.integrity),
      .core_xsecure_ctrl_cpuctrl_pc_hardening                                                                           (core_i.xsecure_ctrl.cpuctrl.pc_hardening),
      .core_xsecure_ctrl_cpuctrl_rndhint                                                                                (core_i.xsecure_ctrl.cpuctrl.rndhint),

      .core_xsecure_ctrl_cpuctrl_rnddummyfreq                                                                           (core_i.xsecure_ctrl.cpuctrl[19:16]),
      .core_if_stage_gen_dummy_instr_dummy_instr_dummy_en                                                               (core_i.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_en),
      .core_cs_registers_xsecure_lfsr_lockup                                                                            (core_i.cs_registers_i.xsecure.lfsr_lockup),

      .core_cs_registers_mhpmcounter_mcycle                                                                             (core_i.cs_registers_i.mcycle_o),
      .core_cs_registers_mhpmcounter_minstret                                                                           (core_i.cs_registers_i.mhpmcounter_q[2]),
      .core_cs_registers_mhpmcounter_31_to_3                                                                            (core_i.cs_registers_i.mhpmcounter_q[31:3]),
      .core_cs_registers_mhpmevent_31_to_3                                                                              (core_i.cs_registers_i.mhpmevent_q[31:3]),
      .core_cs_registers_mcountinhibit_q_mcycle_inhibit                                                                 (core_i.cs_registers_i.mcountinhibit_q[0]),
      .core_cs_registers_mcountinhibit_q_minstret_inhibit                                                               (core_i.cs_registers_i.mcountinhibit_q[2]),

      .core_cs_registers_csr_en_gated                                                                                   (core_i.cs_registers_i.csr_en_gated),
      .core_cs_registers_csr_waddr                                                                                      (core_i.cs_registers_i.csr_waddr),

      .core_LFSR0_CFG_default_seed                                                                                      (core_i.LFSR0_CFG.default_seed),
      .core_LFSR1_CFG_default_seed                                                                                      (core_i.LFSR1_CFG.default_seed),
      .core_LFSR2_CFG_default_seed                                                                                      (core_i.LFSR2_CFG.default_seed),

      .core_xsecure_ctrl_lfsr0                                                                                          (core_i.xsecure_ctrl.lfsr0),
      .core_xsecure_ctrl_lfsr1                                                                                          (core_i.xsecure_ctrl.lfsr1),
      .core_xsecure_ctrl_lfsr2                                                                                          (core_i.xsecure_ctrl.lfsr2),

      .core_cs_registers_xsecure_lfsr0_seed_we                                                                          (core_i.cs_registers_i.xsecure.lfsr0_i.seed_we_i),
      .core_cs_registers_xsecure_lfsr1_seed_we                                                                          (core_i.cs_registers_i.xsecure.lfsr1_i.seed_we_i),
      .core_cs_registers_xsecure_lfsr2_seed_we                                                                          (core_i.cs_registers_i.xsecure.lfsr2_i.seed_we_i),

      .core_i_cs_registers_i_mepc_o                                                                                     (core_i.cs_registers_i.mepc_o),

      // Hardend CSR registers
      .core_i_cs_registers_i_mstateen0_q                                                                                (core_i.cs_registers_i.mstateen0_q),
      .core_i_cs_registers_i_priv_lvl_q_int                                                                             (core_i.cs_registers_i.priv_lvl_q_int),
      .core_i_cs_registers_i_jvt_q                                                                                      (core_i.cs_registers_i.jvt_q),
      .core_i_cs_registers_i_mstatus_q                                                                                  (core_i.cs_registers_i.mstatus_q),
      .core_i_cs_registers_i_cpuctrl_q                                                                                  (core_i.cs_registers_i.cpuctrl_q),
      .core_i_cs_registers_i_dcsr_q                                                                                     (core_i.cs_registers_i.dcsr_q),
      .core_i_cs_registers_i_mepc_q                                                                                     (core_i.cs_registers_i.mepc_q),
      .core_i_cs_registers_i_mscratch_q                                                                                 (core_i.cs_registers_i.mscratch_q),

      .core_i_cs_registers_i_pmp_mseccfg_q                                                                              (core_i.cs_registers_i.pmp_mseccfg_q),
      .core_i_cs_registers_i_pmpncfg_q                                                                                  (core_i.cs_registers_i.pmpncfg_q),
      .core_i_cs_registers_i_pmp_addr_q                                                                                 (core_i.cs_registers_i.pmp_addr_q),

      .core_i_cs_registers_i_mtvt_q                                                                                     (core_i.cs_registers_i.mtvt_q),
      .core_i_cs_registers_i_mtvec_q                                                                                    (core_i.cs_registers_i.mtvec_q),
      .core_i_cs_registers_i_mintstatus_q                                                                               (core_i.cs_registers_i.mintstatus_q),
      .core_i_cs_registers_i_mintthresh_q                                                                               (core_i.cs_registers_i.mintthresh_q),
      .core_i_cs_registers_i_mie_q                                                                                      (core_i.cs_registers_i.mie_q),

      // Shadow registers
      .core_cs_registers_mstateen0_csr_gen_hardened_shadow_q                                                            (core_i.cs_registers_i.mstateen0_csr_i.gen_hardened.shadow_q),
      .core_cs_registers_priv_lvl_gen_hardened_shadow_q                                                                 (core_i.cs_registers_i.priv_lvl_i.gen_hardened.shadow_q),
      .core_cs_registers_jvt_csr_gen_hardened_shadow_q                                                                  (core_i.cs_registers_i.jvt_csr_i.gen_hardened.shadow_q),
      .core_cs_registers_mstatus_csr_gen_hardened_shadow_q                                                              (core_i.cs_registers_i.mstatus_csr_i.gen_hardened.shadow_q),
      .core_cs_registers_xsecure_cpuctrl_csr_gen_hardened_shadow_q                                                      (core_i.cs_registers_i.xsecure.cpuctrl_csr_i.gen_hardened.shadow_q),
      .core_cs_registers_dcsr_csr_gen_hardened_shadow_q                                                                 (core_i.cs_registers_i.dcsr_csr_i.gen_hardened.shadow_q),
      .core_cs_registers_mepc_csr_gen_hardened_shadow_q                                                                 (core_i.cs_registers_i.mepc_csr_i.gen_hardened.shadow_q),
      .core_cs_registers_mscratch_csr_gen_hardened_shadow_q                                                             (core_i.cs_registers_i.mscratch_csr_i.gen_hardened.shadow_q),

      .uvmt_cv32e40s_tb_pmp_mseccfg_q_shadow_q                                                                          (uvmt_cv32e40s_tb.pmp_mseccfg_q_shadow_q),
      .uvmt_cv32e40s_tb_pmpncfg_q_shadow_q                                                                              (uvmt_cv32e40s_tb.pmpncfg_q_shadow_q),
      .uvmt_cv32e40s_tb_pmp_addr_q_shadow_q                                                                             (uvmt_cv32e40s_tb.pmp_addr_q_shadow_q),

      .uvmt_cv32e40s_tb_mtvt_q_shadow_q                                                                                 (uvmt_cv32e40s_tb.mtvt_q_shadow_q),
      .uvmt_cv32e40s_tb_mtvec_q_shadow_q                                                                                (uvmt_cv32e40s_tb.mtvec_q_shadow_q),
      .uvmt_cv32e40s_tb_mintstatus_q_shadow_q                                                                           (uvmt_cv32e40s_tb.mintstatus_q_shadow_q),
      .uvmt_cv32e40s_tb_mintthresh_q_shadow_q                                                                           (uvmt_cv32e40s_tb.mintthresh_q_shadow_q),
      .uvmt_cv32e40s_tb_mie_q_hardened_shadow_q                                                                         (uvmt_cv32e40s_tb.mie_q_hardened_shadow_q),

      // Controller
      .core_i_controller_i_controller_fsm_i_pending_nmi                                                                 (core_i.controller_i.controller_fsm_i.pending_nmi),
      .core_i_controller_i_controller_fsm_i_dcsr_i_step                                                                 (core_i.controller_i.controller_fsm_i.dcsr_i.step),
      .core_i_controller_i_controller_fsm_i_dcsr_i_stepie                                                                 (core_i.controller_i.controller_fsm_i.dcsr_i.stepie),
      .core_controller_controller_fsm_debug_mode_q                                                                      (core_i.controller_i.controller_fsm_i.debug_mode_q),

      // IF stage
      .core_if_stage_if_valid_o                                                                                         (core_i.if_stage_i.if_valid_o),
      .core_if_stage_id_ready_i                                                                                         (core_i.if_stage_i.id_ready_i),

      .core_if_stage_gen_dummy_instr_dummy_instr_lfsr_rs1                                                               (core_i.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_rs1),
      .core_if_stage_gen_dummy_instr_dummy_instr_lfsr_rs2                                                               (core_i.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_rs2),

      .core_if_stage_instr_meta_n_dummy                                                                                 (core_i.if_stage_i.instr_meta_n.dummy),
      .core_i_if_stage_i_instr_hint                                                                                     (core_i.if_stage_i.instr_hint),
      .core_i_if_stage_i_dummy_insert                                                                                   (core_i.if_stage_i.dummy_insert),

      .core_i_if_stage_i_pc_if_o                                                                                        (core_i.if_stage_i.pc_if_o),
      .core_i_if_stage_i_pc_check_i_pc_set_q                                                                            (core_i.if_stage_i.pc_check_i.pc_set_q),

      .core_i_if_stage_i_ptr_in_if_o                                                                                    (core_i.if_stage_i.ptr_in_if_o),
      .core_i_if_stage_i_compressed_decoder_i_is_compressed_o                                                           (core_i.if_stage_i.compressed_decoder_i.is_compressed_o),

      // IF ID pipe
      .core_if_id_pipe_instr_meta_dummy                                                                                 (core_i.if_id_pipe.instr_meta.dummy),
      .core_if_id_pipe_instr_meta_hint                                                                                  (core_i.if_id_pipe.instr_meta.hint),
      .core_if_id_pipe_instr_bus_resp_rdata                                                                             (core_i.if_id_pipe.instr.bus_resp.rdata),
      .core_i_id_stage_i_if_id_pipe_i_pc                                                                                (core_i.id_stage_i.if_id_pipe_i.pc),
      .core_i_if_id_pipe_last_op                                                                                        (core_i.if_id_pipe.last_op),

      // ID stage
      .core_id_stage_id_valid_o                                                                                         (core_i.id_stage_i.id_valid_o),
      .core_id_stage_ex_ready_i                                                                                         (core_i.id_stage_i.ex_ready_i),
      .core_id_stage_if_id_pipe_instr_meta_compressed                                                                   (core_i.id_stage_i.if_id_pipe_i.instr_meta.compressed),
      .core_id_stage_if_id_pipe_compressed_instr                                                                        (core_i.id_stage_i.if_id_pipe_i.compressed_instr),

      // ID EX pipe
      .core_id_ex_pipe_instr_meta_dummy                                                                                 (core_i.id_ex_pipe.instr_meta.dummy),

      // EX stage
      .core_i_ex_stage_i_branch_target_o                                                                                (core_i.ex_stage_i.branch_target_o),
      .core_i_ex_stage_i_alu_i_cmp_result_o                                                                             (core_i.ex_stage_i.alu_i.cmp_result_o),

      // EX WB pipe
      .core_ex_wb_pipe_instr_meta_dummy                                                                                 (core_i.ex_wb_pipe.instr_meta.dummy),
      .core_ex_wb_pipe_instr_meta_hint                                                                                  (core_i.ex_wb_pipe.instr_meta.hint),

      // WB stage
      .core_wb_stage_wb_valid_o                                                                                         (core_i.wb_stage_i.wb_valid_o),

      // CTRL
      .core_i_if_stage_i_prefetch_unit_i_alignment_buffer_i_ctrl_fsm_i_pc_set                                           (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.ctrl_fsm_i.pc_set),
      .core_i_if_stage_i_pc_check_i_ctrl_fsm_i_pc_mux                                                                   (core_i.if_stage_i.pc_check_i.ctrl_fsm_i.pc_mux)

    );
   // Xsecure assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_xsecure_assert #(
      .SECURE              (cv32e40s_pkg::SECURE),
      .SMCLIC              (SMCLIC),
      .PMP_NUM_REGIONS     (PMP_NUM_REGIONS),
      .MTVT_ADDR_WIDTH     (core_i.MTVT_ADDR_WIDTH),
      .CSR_MINTTHRESH_MASK (core_i.cs_registers_i.CSR_MINTTHRESH_MASK),
      .PMP_ADDR_WIDTH      (core_i.cs_registers_i.PMP_ADDR_WIDTH)
    ) xsecure_assert_i (
      .clk_i      (clknrst_if.clk),
      .rst_ni     (clknrst_if.reset_n),
      .xsecure_if (xsecure_if),
      .rvfi_if    (rvfi_instr_if_0_i),
      .support_if (support_logic_for_assert_coverage_modules_if.slave_mp)
    );

  // Debug assertion and coverage interface

  // Instantiate debug assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_debug_cov_assert_if  debug_cov_assert_if (
      .id_valid               (core_i.id_stage_i.id_valid_o),
      .sys_fence_insn_i       (core_i.id_stage_i.decoder_i.sys_fencei_insn_o),

      .ex_stage_csr_en        (core_i.id_ex_pipe.csr_en),
      .ex_valid               (core_i.ex_stage_i.instr_valid),
      .ex_stage_instr_rdata_i (core_i.id_ex_pipe.instr.bus_resp.rdata),
      .ex_stage_pc            (core_i.id_ex_pipe.pc),

      .wb_stage_instr_rdata_i (core_i.ex_wb_pipe.instr.bus_resp.rdata),
      .wb_stage_instr_valid_i (core_i.ex_wb_pipe.instr_valid),
      .wb_stage_pc            (core_i.wb_stage_i.ex_wb_pipe_i.pc),
      .wb_err                 (core_i.ex_wb_pipe.instr.bus_resp.err),
      .wb_illegal             (core_i.ex_wb_pipe.illegal_insn),
      .wb_valid               (core_i.wb_stage_i.wb_valid_o),
      .wb_mpu_status          (core_i.ex_wb_pipe.instr.mpu_status),
      .illegal_insn_i         (core_i.ex_wb_pipe.illegal_insn),
      .sys_en_i               (core_i.ex_wb_pipe.sys_en),
      .sys_ecall_insn_i       (core_i.ex_wb_pipe.sys_ecall_insn),

      .ctrl_fsm_cs            (core_i.controller_i.controller_fsm_i.ctrl_fsm_cs),
      .debug_req_i            (core_i.controller_i.controller_fsm_i.debug_req_i),
      .debug_havereset        (core_i.debug_havereset_o),
      .debug_running          (core_i.debug_running_o),
      .debug_halted           (core_i.debug_halted_o),

      .ctrl_fsm_async_debug_allowed  (core_i.controller_i.controller_fsm_i.async_debug_allowed),
      .pending_sync_debug     (core_i.controller_i.controller_fsm_i.pending_sync_debug),
      .pending_async_debug    (core_i.controller_i.controller_fsm_i.pending_async_debug),
      .pending_nmi            (core_i.controller_i.controller_fsm_i.pending_nmi),
      .nmi_allowed            (core_i.controller_i.controller_fsm_i.nmi_allowed),
      .debug_mode_q           (core_i.controller_i.controller_fsm_i.debug_mode_q),
      .trigger_match_in_wb    (core_i.controller_i.controller_fsm_i.trigger_match_in_wb),
      .etrigger_in_wb         (core_i.controller_i.controller_fsm_i.etrigger_in_wb),
      .branch_in_ex           (core_i.controller_i.controller_fsm_i.branch_in_ex),

      .mie_q                  (core_i.cs_registers_i.mie_q),
      .dcsr_q                 (core_i.cs_registers_i.dcsr_q),
      .dpc_q                  (core_i.cs_registers_i.dpc_q),
      .dpc_n                  (core_i.cs_registers_i.dpc_n),
      .mcause_q               (core_i.cs_registers_i.mcause_q),
      .mtvec                  (core_i.cs_registers_i.mtvec_q),
      .mepc_q                 (core_i.cs_registers_i.mepc_q),
      .tdata1                 (core_i.cs_registers_i.tdata1_rdata),
      .tdata2                 (core_i.cs_registers_i.tdata2_rdata),
      .mcountinhibit_q        (core_i.cs_registers_i.mcountinhibit_q),
      .mcycle                 (core_i.cs_registers_i.mhpmcounter_q[0]),
      .minstret               (core_i.cs_registers_i.mhpmcounter_q[2]),
      .csr_we_int             (core_i.cs_registers_i.csr_we_int),

      // TODO: review this change from CV32E40S_HASH f6196bf to a26b194. It should be logically equivalent.
      //assign debug_cov_assert_if.inst_ret = core_i.cs_registers_i.inst_ret;
      // First attempt: this causes unexpected failures of a_minstret_count
      //assign debug_cov_assert_if.inst_ret = (core_i.id_valid &
      //                                       core_i.is_decoding);
      // Second attempt: (based on OK input).  This passes, but maybe only because p_minstret_count
      //                                       is the only property sensitive to inst_ret. Will
      //                                       this work in the general case?
      .inst_ret               (core_i.ctrl_fsm.mhpmevent.minstret),
      .csr_access             (core_i.ex_wb_pipe.csr_en),
      .csr_op                 (core_i.ex_wb_pipe.csr_op),
      .csr_addr               (core_i.ex_wb_pipe.csr_addr),
      .irq_ack_o              (core_i.irq_ack),
      .irq_id_o               (core_i.irq_id),
      .dm_halt_addr_i         (core_i.dm_halt_addr_i),
      .dm_exception_addr_i    (core_i.dm_exception_addr_i),
      .core_sleep_o           (core_i.core_sleep_o),
      .irq_i                  (core_i.irq_i),
      .pc_set                 (core_i.ctrl_fsm.pc_set),
      .boot_addr_i            (core_i.boot_addr_i),

      .is_wfi                 (),
      .dpc_will_hit           (),
      .addr_match             (),
      .is_ebreak              (),
      .is_cebreak             (),
      .is_dret                (),
      .is_mulhsu              (),
      .pending_enabled_irq    (),

      .*
    );


    bind cv32e40s_wrapper
      uvmt_cv32e40s_input_to_support_logic_module_if input_to_support_logic_module_if (
        .clk     (core_i.clk),
        .rst_n (rst_ni),

        .ctrl_fsm_o (core_i.controller_i.controller_fsm_i.ctrl_fsm_o),

        .data_bus_rvalid (core_i.m_c_obi_data_if.s_rvalid.rvalid),
        .data_bus_req (core_i.m_c_obi_data_if.s_req.req),
        .data_bus_gnt (core_i.m_c_obi_data_if.s_gnt.gnt),
        .data_bus_gntpar (core_i.m_c_obi_data_if.s_gnt.gntpar),

        .instr_bus_rvalid (core_i.m_c_obi_instr_if.s_rvalid.rvalid),
        .instr_bus_req (core_i.m_c_obi_instr_if.s_req.req),
        .instr_bus_gnt (core_i.m_c_obi_instr_if.s_gnt.gnt),
        .instr_bus_gntpar (core_i.m_c_obi_instr_if.s_gnt.gntpar),

        //obi protocol between alignmentbuffer (ab) and instructoin (i) interface (i) mpu (m) is refered to as abiim
        .abiim_bus_rvalid (core_i.if_stage_i.prefetch_resp_valid),
        .abiim_bus_req (core_i.if_stage_i.prefetch_trans_ready),
        .abiim_bus_gnt (core_i.if_stage_i.prefetch_trans_valid),

        //obi protocol between LSU (l) mpu (m) and LSU (l) is refered to as lml
        .lml_bus_rvalid (core_i.load_store_unit_i.resp_valid),
        .lml_bus_req (core_i.load_store_unit_i.trans_ready),
        .lml_bus_gnt (core_i.load_store_unit_i.trans_valid),

        //obi protocol between LSU (l) respons (r) filter (f) and OBI (o) data (d) interface (i) is refered to as lrfodi
        .lrfodi_bus_rvalid (core_i.load_store_unit_i.bus_resp_valid),
        .lrfodi_bus_req (core_i.load_store_unit_i.buffer_trans_valid),
        .lrfodi_bus_gnt (core_i.load_store_unit_i.buffer_trans_ready),

        .req_is_store (core_i.load_store_unit_i.bus_trans.we),
        .req_instr_integrity (core_i.if_stage_i.mpu_i.bus_trans_integrity),
        .req_data_integrity (core_i.load_store_unit_i.mpu_i.bus_trans_integrity)

    );

    bind cv32e40s_wrapper
      uvmt_cv32e40s_support_logic_for_assert_coverage_modules_if support_logic_for_assert_coverage_modules_if();

    bind cv32e40s_pmp :
      uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i.pmp.pmp_i
      uvmt_cv32e40s_pmp_assert #(
        .PMP_GRANULARITY  (PMP_GRANULARITY),
        .PMP_NUM_REGIONS  (PMP_NUM_REGIONS),
        .IS_INSTR_SIDE    (1'b1),
        .PMP_MSECCFG_RV   (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_MSECCFG_RV)
      )
      u_pmp_assert_if_stage(.rst_n          (clknrst_if.reset_n),
                            .bus_trans_dbg  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i.bus_trans_o.dbg),
                            .obi_addr       (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_addr_o),
                            .obi_gnt        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_gnt_i),
                            .obi_req        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_req_o),
                            .rvfi_pc_rdata  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_pc_rdata),
                            .rvfi_valid     (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_valid),
                            .*);

    bind  cv32e40s_pmp :
      uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i.pmp.pmp_i
      uvmt_cv32e40s_pmp_assert#(
        .PMP_GRANULARITY  (PMP_GRANULARITY),
        .PMP_NUM_REGIONS  (PMP_NUM_REGIONS),
        .IS_INSTR_SIDE    (1'b0),
        .PMP_MSECCFG_RV   (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_MSECCFG_RV)
      )
      u_pmp_assert_lsu(.rst_n          (clknrst_if.reset_n),
                       .bus_trans_dbg  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i.bus_trans_o.dbg),
                       .obi_addr       (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_addr_o),
                       .obi_gnt        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_gnt_i),
                       .obi_req        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_req_o),
                       .rvfi_pc_rdata  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_pc_rdata),
                       .rvfi_valid     (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_valid),
                       .*);

    bind  dut_wrap.cv32e40s_wrapper_i.rvfi_i
      uvmt_cv32e40s_pmprvfi_assert #(
        .PMP_GRANULARITY (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_GRANULARITY),
        .PMP_NUM_REGIONS (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_NUM_REGIONS)
      ) pmprvfi_assert_i (
        .rvfi_mem_addr  (rvfi_mem_addr [31:0]),
        .rvfi_mem_wmask (rvfi_mem_wmask[ 3:0]),
        .rvfi_mem_rmask (rvfi_mem_rmask[ 3:0]),
        .*
      );

    bind  dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i
      uvmt_cv32e40s_pma_assert #(
        .CORE_REQ_TYPE   (cv32e40s_pkg::obi_inst_req_t),
        .DM_REGION_END   (uvmt_cv32e40s_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (1),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_CFG)
      ) pma_assert_instr_i (
        .obi              (dut_wrap.obi_instr_if_i),
        .rvfi             (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i),
        .sup              (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.support_logic_for_assert_coverage_modules_if),
        .writebuf_ready_o ('0),
        .writebuf_trans_i ('0),
        .writebuf_trans_o ('0),
        .*
      );

    bind  dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i
      uvmt_cv32e40s_pma_assert #(
        .CORE_REQ_TYPE   (cv32e40s_pkg::obi_data_req_t),
        .DM_REGION_END   (uvmt_cv32e40s_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (0),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_CFG)
      ) pma_assert_data_i (
        .obi              (dut_wrap.obi_data_if_i),
        .rvfi             (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i),
        .sup              (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.support_logic_for_assert_coverage_modules_if),
        .writebuf_ready_o (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.ready_o),
        .writebuf_trans_i (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.trans_i),
        .writebuf_trans_o (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.trans_o),
        .*
      );

    bind cv32e40s_wrapper uvmt_cv32e40s_support_logic u_support_logic(.rvfi(rvfi_instr_if_0_i),
                                                                      .in_support_if (input_to_support_logic_module_if.driver_mp),
                                                                      .out_support_if (support_logic_for_assert_coverage_modules_if.master_mp)
                                                                      );

    bind cv32e40s_wrapper uvmt_cv32e40s_debug_assert u_debug_assert(.rvfi(rvfi_instr_if_0_i),
                                                                    .csr_dcsr(rvfi_csr_dcsr_if_0_i),
                                                                    .csr_dpc(rvfi_csr_dpc_if_0_i),
                                                                    .csr_mepc(rvfi_csr_mepc_if_0_i),
                                                                    .csr_mstatus(rvfi_csr_mstatus_if_0_i),
                                                                    .csr_mtvec(rvfi_csr_mtvec_if_0_i),
                                                                    .csr_tdata1(rvfi_csr_tdata1_if_0_i),
                                                                    .cov_assert_if(debug_cov_assert_if));

    bind cv32e40s_wrapper uvmt_cv32e40s_zc_assert u_zc_assert(.rvfi(rvfi_instr_if_0_i),
                                                              .support_if(support_logic_for_assert_coverage_modules_if.slave_mp)
                                                              );


    //uvmt_cv32e40s_rvvi_handcar u_rvvi_handcar();

    // IMPERAS DV
    `ifndef FORMAL
      uvmt_cv32e40s_imperas_dv_wrap imperas_dv (rvvi_if);
    `endif

   /**
    * Test bench entry point.
    */
   `ifndef FORMAL // Formal ignores initial blocks, avoids unnecessary warning
   initial begin : test_bench_entry_point

     // Specify time format for simulation (units_number, precision_number, suffix_string, minimum_field_width)
     $timeformat(-9, 3, " ns", 8);

     // Add interfaces handles to uvm_config_db
     uvm_config_db#(virtual uvma_isacov_if              )::set(.cntxt(null), .inst_name("*.env.isacov_agent"),           .field_name("vif"),           .value(isacov_if));
     uvm_config_db#(virtual uvma_debug_if               )::set(.cntxt(null), .inst_name("*.env.debug_agent"),            .field_name("vif"),           .value(debug_if));
     uvm_config_db#(virtual uvma_clknrst_if             )::set(.cntxt(null), .inst_name("*.env.clknrst_agent"),          .field_name("vif"),           .value(clknrst_if));
     uvm_config_db#(virtual uvma_interrupt_if           )::set(.cntxt(null), .inst_name("*.env.interrupt_agent"),        .field_name("vif"),           .value(interrupt_if));
     uvm_config_db#(virtual uvma_clic_if                )::set(.cntxt(null), .inst_name("*.env.clic_agent"),             .field_name("vif"),           .value(clic_if));

     uvm_config_db#(virtual uvma_obi_memory_if#(
       .AUSER_WIDTH(ENV_PARAM_INSTR_AUSER_WIDTH),
       .WUSER_WIDTH(ENV_PARAM_INSTR_WUSER_WIDTH),
       .RUSER_WIDTH(ENV_PARAM_INSTR_RUSER_WIDTH),
       .ADDR_WIDTH(ENV_PARAM_INSTR_ADDR_WIDTH),
       .DATA_WIDTH(ENV_PARAM_INSTR_DATA_WIDTH),
       .ID_WIDTH(ENV_PARAM_INSTR_ID_WIDTH),
       .ACHK_WIDTH(ENV_PARAM_INSTR_ACHK_WIDTH),
       .RCHK_WIDTH(ENV_PARAM_INSTR_RCHK_WIDTH)
     ))::set(.cntxt(null), .inst_name("*.env.obi_memory_instr_agent"), .field_name("vif"), .value(obi_instr_if_i) );
     uvm_config_db#(virtual uvma_obi_memory_if#(
       .AUSER_WIDTH(ENV_PARAM_DATA_AUSER_WIDTH),
       .WUSER_WIDTH(ENV_PARAM_DATA_WUSER_WIDTH),
       .RUSER_WIDTH(ENV_PARAM_DATA_RUSER_WIDTH),
       .ADDR_WIDTH(ENV_PARAM_DATA_ADDR_WIDTH),
       .DATA_WIDTH(ENV_PARAM_DATA_DATA_WIDTH),
       .ID_WIDTH(ENV_PARAM_DATA_ID_WIDTH),
       .ACHK_WIDTH(ENV_PARAM_DATA_ACHK_WIDTH),
       .RCHK_WIDTH(ENV_PARAM_DATA_RCHK_WIDTH)
     ))::set(.cntxt(null), .inst_name("*.env.obi_memory_data_agent"),  .field_name("vif"), .value(obi_data_if_i) );
     uvm_config_db#(virtual uvma_fencei_if              )::set(.cntxt(null), .inst_name("*.env.fencei"),                 .field_name("vif"),           .value(fencei_if_i));
     uvm_config_db#(virtual uvma_rvfi_instr_if          )::set(.cntxt(null), .inst_name("*.env.rvfi_agent"),             .field_name("instr_vif0"),    .value(dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i));
     uvm_config_db#(virtual uvma_fencei_if              )::set(.cntxt(null), .inst_name("*.env.fencei_agent"),           .field_name("fencei_vif"),    .value(fencei_if_i)  );
     uvm_config_db#(virtual uvmt_cv32e40s_vp_status_if  )::set(.cntxt(null), .inst_name("*"),                            .field_name("vp_status_vif"), .value(vp_status_if) );
     uvm_config_db#(virtual uvma_interrupt_if           )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("intr_vif"),      .value(interrupt_if) );
     uvm_config_db#(virtual uvma_clic_if                )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("clic_vif"),      .value(clic_if) );
     uvm_config_db#(virtual uvma_debug_if               )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("debug_vif"),     .value(debug_if)     );
//     uvm_config_db#(virtual uvmt_cv32e40s_debug_cov_assert_if)::set(.cntxt(null), .inst_name("*.env"),                 .field_name("debug_cov_vif"),    .value(debug_cov_assert_if));
     `RVFI_CSR_UVM_CONFIG_DB_SET(cpuctrl)
     `RVFI_CSR_UVM_CONFIG_DB_SET(jvt)
     `RVFI_CSR_UVM_CONFIG_DB_SET(marchid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcause)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcounteren)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcountinhibit)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcycle)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcycleh)
     `RVFI_CSR_UVM_CONFIG_DB_SET(menvcfg)
     `RVFI_CSR_UVM_CONFIG_DB_SET(menvcfgh)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mepc)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhartid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mie)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mimpid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(minstret)
     `RVFI_CSR_UVM_CONFIG_DB_SET(minstreth)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mip)
     `RVFI_CSR_UVM_CONFIG_DB_SET(misa)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mscratch)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen0h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen1h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen2h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen3h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstatus)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstatush)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mtval)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mtvec)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mvendorid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mseccfg)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mseccfgh)

     `RVFI_CSR_UVM_CONFIG_DB_SET(dcsr)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dpc)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dscratch0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dscratch1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tselect)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tinfo)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tcontrol)

     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg15)

     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr31)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr32)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr33)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr34)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr35)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr36)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr37)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr38)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr39)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr40)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr41)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr42)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr43)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr44)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr45)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr46)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr47)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr48)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr49)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr50)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr51)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr52)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr53)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr54)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr55)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr56)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr57)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr58)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr59)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr60)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr61)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr62)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr63)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent31)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter31)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter3h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter4h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter5h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter6h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter7h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter8h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter9h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter10h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter11h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter12h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter13h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter14h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter15h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter16h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter17h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter18h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter19h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter20h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter21h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter22h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter23h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter24h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter25h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter26h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter27h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter28h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter29h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter30h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter31h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mconfigptr)

     `RVFI_CSR_UVM_CONFIG_DB_SET(secureseed0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(secureseed1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(secureseed2)

     `ifdef SMCLIC_EN
       // TODO:silabs-robin  What about when using "PARAM_SET_0"?
       `RVFI_CSR_UVM_CONFIG_DB_SET(mintstatus)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mintthresh)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mnxti)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mscratchcsw)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mscratchcswl)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mtvt)
     `endif

     // IMPERAS_DV interface
     uvm_config_db#(virtual rvviTrace)::set(.cntxt(null), .inst_name("*.env.rvvi_agent"), .field_name("rvvi_vif"), .value(rvvi_if));

     // Virtual Peripheral Status interface
     uvm_config_db#(virtual uvmt_cv32e40s_vp_status_if      )::set(.cntxt(null), .inst_name("*"), .field_name("vp_status_vif"),       .value(vp_status_if)      );
     uvm_config_db#(virtual uvme_cv32e40s_core_cntrl_if     )::set(.cntxt(null), .inst_name("*"), .field_name("core_cntrl_vif"),      .value(core_cntrl_if)     );
     uvm_config_db#(virtual uvmt_cv32e40s_core_status_if    )::set(.cntxt(null), .inst_name("*"), .field_name("core_status_vif"),     .value(core_status_if)    );
     uvm_config_db#(virtual uvmt_cv32e40s_debug_cov_assert_if)::set(.cntxt(null), .inst_name("*.env"), .field_name("debug_cov_vif"),.value(dut_wrap.cv32e40s_wrapper_i.debug_cov_assert_if));
     uvm_config_db#(virtual uvmt_cv32e40s_support_logic_for_assert_coverage_modules_if)::set(.cntxt(null), .inst_name("*.env"), .field_name("support_logic_vif"),.value(dut_wrap.cv32e40s_wrapper_i.support_logic_for_assert_coverage_modules_if));

     // Make the DUT Wrapper Virtual Peripheral's status outputs available to the base_test
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("tp"),     .value(1'b0)        );
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("tf"),     .value(1'b0)        );
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("evalid"), .value(1'b0)        );
     uvm_config_db#(bit[31:0])::set(.cntxt(null), .inst_name("*"), .field_name("evalue"), .value(32'h00000000));

	   // DUT and ENV parameters
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_INSTR_ADDR_WIDTH"),  .value(ENV_PARAM_INSTR_ADDR_WIDTH) );
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_INSTR_DATA_WIDTH"),  .value(ENV_PARAM_INSTR_DATA_WIDTH) );
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_RAM_ADDR_WIDTH"),    .value(ENV_PARAM_RAM_ADDR_WIDTH)   );

     // Run test
     uvm_top.enable_print_topology = 0; // ENV coders enable this as a debug aid
     uvm_top.finish_on_completion  = 1;
     uvm_top.run_test();
   end : test_bench_entry_point
   `endif

   assign core_cntrl_if.clk = clknrst_if.clk;

   // Informational print message on loading of OVPSIM ISS to benchmark some elf image loading times
   // OVPSIM runs its initialization at the #1ns timestamp, and should dominate the initial startup time
   `ifndef FORMAL // Formal ignores initial blocks, avoids unnecessary warning
   // overcome race
   initial begin
     if ($test$plusargs("USE_ISS")) begin
       #0.9ns;
       imperas_dv.ref_init();
     end
   end
   `endif

   //TODO verify these are correct with regards to isacov function
   `ifndef FORMAL // events ignored for formal - this avoids unnecessary warning
     always @(dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i.rvfi_valid) -> isacov_if.retire;
   `endif
   assign isacov_if.instr = dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i.rvfi_insn;
   //assign isacov_if.is_compressed = dut_wrap.cv32e40s_wrapper_i.tracer_i.insn_compressed;

   // Capture the test status and exit pulse flags
   // TODO: put this logic in the vp_status_if (makes it easier to pass to ENV)
   `ifndef FORMAL  // uvm db not used in formal
     always @(posedge clknrst_if.clk) begin
       if (!clknrst_if.reset_n) begin
         tp     <= 1'b0;
         tf     <= 1'b0;
         evalid <= 1'b0;
         evalue <= 32'h00000000;
       end
       else begin
         if (vp_status_if.tests_passed) begin
           tp <= 1'b1;
           uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("tp"), .value(1'b1));
         end
         if (vp_status_if.tests_failed) begin
           tf <= 1'b1;
           uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("tf"), .value(1'b1));
         end
         if (vp_status_if.exit_valid) begin
           evalid <= 1'b1;
           uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("evalid"), .value(1'b1));
         end
         if (vp_status_if.exit_valid) begin
           evalue <= vp_status_if.exit_value;
           uvm_config_db#(bit[31:0])::set(.cntxt(null), .inst_name("*"), .field_name("evalue"), .value(vp_status_if.exit_value));
         end
       end
     end
   `endif  // FORMAL


   /**
    * End-of-test summary printout.
    */
   `ifndef FORMAL // Formal ignores final blocks, this avoids unnecessary warning
   final begin: end_of_test
      string             summary_string;
      uvm_report_server  rs;
      int                err_count;
      int                warning_count;
      int                fatal_count;
      static bit         sim_finished = 0;

      static string  red   = "\033[31m\033[1m";
      static string  green = "\033[32m\033[1m";
      static string  reset = "\033[0m";

      rs            = uvm_top.get_report_server();
      err_count     = rs.get_severity_count(UVM_ERROR);
      warning_count = rs.get_severity_count(UVM_WARNING);
      fatal_count   = rs.get_severity_count(UVM_FATAL);

      void'(uvm_config_db#(bit)::get(null, "", "sim_finished", sim_finished));

      // Shutdown the Reference Model
      if ($test$plusargs("USE_ISS")) begin
         // Exit handler for ImperasDV
         void'(rvviRefShutdown());
      end

      `uvm_info("DV_WRAP", $sformatf("\n%m: *** Test Summary ***\n"), UVM_DEBUG);

      if (sim_finished && (err_count == 0) && (fatal_count == 0)) begin
         $display("    PPPPPPP    AAAAAA    SSSSSS    SSSSSS   EEEEEEEE  DDDDDDD     ");
         $display("    PP    PP  AA    AA  SS    SS  SS    SS  EE        DD    DD    ");
         $display("    PP    PP  AA    AA  SS        SS        EE        DD    DD    ");
         $display("    PPPPPPP   AAAAAAAA   SSSSSS    SSSSSS   EEEEE     DD    DD    ");
         $display("    PP        AA    AA        SS        SS  EE        DD    DD    ");
         $display("    PP        AA    AA  SS    SS  SS    SS  EE        DD    DD    ");
         $display("    PP        AA    AA   SSSSSS    SSSSSS   EEEEEEEE  DDDDDDD     ");
         $display("    ----------------------------------------------------------");
         if (warning_count == 0) begin
           $display("                        SIMULATION PASSED                     ");
         end
         else begin
           $display("                 SIMULATION PASSED with WARNINGS              ");
         end
         $display("    ----------------------------------------------------------");
      end
      else begin
         $display("    FFFFFFFF   AAAAAA   IIIIII  LL        EEEEEEEE  DDDDDDD       ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FFFFF     AAAAAAAA    II    LL        EEEEE     DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA  IIIIII  LLLLLLLL  EEEEEEEE  DDDDDDD       ");

         if (sim_finished == 0) begin
            $display("    --------------------------------------------------------");
            $display("                   SIMULATION FAILED - ABORTED              ");
            $display("    --------------------------------------------------------");
         end
         else begin
            $display("    --------------------------------------------------------");
            $display("                       SIMULATION FAILED                    ");
            $display("    --------------------------------------------------------");
         end
      end
   end
   `endif

endmodule : uvmt_cv32e40s_tb
`default_nettype wire

`endif // __UVMT_CV32E40S_TB_SV__
