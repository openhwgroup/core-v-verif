// ----------------------------------------------------------------------------
//Copyright 2023 CEA*
//*Commissariat a l'Energie Atomique et aux Energies Alternatives (CEA)
//
//Licensed under the Apache License, Version 2.0 (the "License");
//you may not use this file except in compliance with the License.
//You may obtain a copy of the License at
//
//    http://www.apache.org/licenses/LICENSE-2.0
//
//Unless required by applicable law or agreed to in writing, software
//distributed under the License is distributed on an "AS IS" BASIS,
//WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//See the License for the specific language governing permissions and
//limitations under the License.
//[END OF HEADER]
// ----------------------------------------------------------------------------
//  Description :
//
//
//  Copyright (C) 2019 CEA-Leti
//  Author      : $authorname : PERBOST Nicolas $ $authoremail : nicolas.perbost.fr $
//
//  Id          : $Id: ebc1c90d292c16718a5f425063aa10baa9553215 $
//  Date        : $Date : Tue Mar 5 17:22:29 2019 +0100 $
//
// ----------------------------------------------------------------------------

package test_pkg;

    import uvm_pkg::*;
    import uvma_axi_pkg::*;
    import dut_env_pkg::*;
    `include "uvm_macros.svh";
    `include "base_test_c.svh";
    `include "bursty_test_c.svh";


endpackage : test_pkg


