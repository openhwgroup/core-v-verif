package uvm_pkg;
endpackage

`define  uvm_error(ID, MSG)  ;
