// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2020 Silicon Labs, Inc.
// Copyright 2023 Thales DIS
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`ifndef __UVMA_CVXIF_MACROS_SV__
`define __UVMA_CVXIF_MACROS_SV__


`define CVXIF_CP_BITWISE_IFF(name, field, iff_exp) \
``name``: coverpoint(``field``) { \
    wildcard bins BIT0_0  = {32'b???????????????????????????????0} with (``iff_exp``); \
    wildcard bins BIT1_0  = {32'b??????????????????????????????0?} with (``iff_exp``); \
    wildcard bins BIT2_0  = {32'b?????????????????????????????0??} with (``iff_exp``); \
    wildcard bins BIT3_0  = {32'b????????????????????????????0???} with (``iff_exp``); \
    wildcard bins BIT4_0  = {32'b???????????????????????????0????} with (``iff_exp``); \
    wildcard bins BIT5_0  = {32'b??????????????????????????0?????} with (``iff_exp``); \
    wildcard bins BIT6_0  = {32'b?????????????????????????0??????} with (``iff_exp``); \
    wildcard bins BIT7_0  = {32'b????????????????????????0???????} with (``iff_exp``); \
    wildcard bins BIT8_0  = {32'b???????????????????????0????????} with (``iff_exp``); \
    wildcard bins BIT9_0  = {32'b??????????????????????0?????????} with (``iff_exp``); \
    wildcard bins BIT10_0 = {32'b?????????????????????0??????????} with (``iff_exp``); \
    wildcard bins BIT11_0 = {32'b????????????????????0???????????} with (``iff_exp``); \
    wildcard bins BIT12_0 = {32'b???????????????????0????????????} with (``iff_exp``); \
    wildcard bins BIT13_0 = {32'b??????????????????0?????????????} with (``iff_exp``); \
    wildcard bins BIT14_0 = {32'b?????????????????0??????????????} with (``iff_exp``); \
    wildcard bins BIT15_0 = {32'b????????????????0???????????????} with (``iff_exp``); \
    wildcard bins BIT16_0 = {32'b???????????????0????????????????} with (``iff_exp``); \
    wildcard bins BIT17_0 = {32'b??????????????0?????????????????} with (``iff_exp``); \
    wildcard bins BIT18_0 = {32'b?????????????0??????????????????} with (``iff_exp``); \
    wildcard bins BIT19_0 = {32'b????????????0???????????????????} with (``iff_exp``); \
    wildcard bins BIT20_0 = {32'b???????????0????????????????????} with (``iff_exp``); \
    wildcard bins BIT21_0 = {32'b??????????0?????????????????????} with (``iff_exp``); \
    wildcard bins BIT22_0 = {32'b?????????0??????????????????????} with (``iff_exp``); \
    wildcard bins BIT23_0 = {32'b????????0???????????????????????} with (``iff_exp``); \
    wildcard bins BIT24_0 = {32'b???????0????????????????????????} with (``iff_exp``); \
    wildcard bins BIT25_0 = {32'b??????0?????????????????????????} with (``iff_exp``); \
    wildcard bins BIT26_0 = {32'b?????0??????????????????????????} with (``iff_exp``); \
    wildcard bins BIT27_0 = {32'b????0???????????????????????????} with (``iff_exp``); \
    wildcard bins BIT28_0 = {32'b???0????????????????????????????} with (``iff_exp``); \
    wildcard bins BIT29_0 = {32'b??0?????????????????????????????} with (``iff_exp``); \
    wildcard bins BIT30_0 = {32'b?0??????????????????????????????} with (``iff_exp``); \
    wildcard bins BIT31_0 = {32'b0???????????????????????????????} with (``iff_exp``); \
    wildcard bins BIT0_1  = {32'b???????????????????????????????1} with (``iff_exp``); \
    wildcard bins BIT1_1  = {32'b??????????????????????????????1?} with (``iff_exp``); \
    wildcard bins BIT2_1  = {32'b?????????????????????????????1??} with (``iff_exp``); \
    wildcard bins BIT3_1  = {32'b????????????????????????????1???} with (``iff_exp``); \
    wildcard bins BIT4_1  = {32'b???????????????????????????1????} with (``iff_exp``); \
    wildcard bins BIT5_1  = {32'b??????????????????????????1?????} with (``iff_exp``); \
    wildcard bins BIT6_1  = {32'b?????????????????????????1??????} with (``iff_exp``); \
    wildcard bins BIT7_1  = {32'b????????????????????????1???????} with (``iff_exp``); \
    wildcard bins BIT8_1  = {32'b???????????????????????1????????} with (``iff_exp``); \
    wildcard bins BIT9_1  = {32'b??????????????????????1?????????} with (``iff_exp``); \
    wildcard bins BIT10_1 = {32'b?????????????????????1??????????} with (``iff_exp``); \
    wildcard bins BIT11_1 = {32'b????????????????????1???????????} with (``iff_exp``); \
    wildcard bins BIT12_1 = {32'b???????????????????1????????????} with (``iff_exp``); \
    wildcard bins BIT13_1 = {32'b??????????????????1?????????????} with (``iff_exp``); \
    wildcard bins BIT14_1 = {32'b?????????????????1??????????????} with (``iff_exp``); \
    wildcard bins BIT15_1 = {32'b????????????????1???????????????} with (``iff_exp``); \
    wildcard bins BIT16_1 = {32'b???????????????1????????????????} with (``iff_exp``); \
    wildcard bins BIT17_1 = {32'b??????????????1?????????????????} with (``iff_exp``); \
    wildcard bins BIT18_1 = {32'b?????????????1??????????????????} with (``iff_exp``); \
    wildcard bins BIT19_1 = {32'b????????????1???????????????????} with (``iff_exp``); \
    wildcard bins BIT20_1 = {32'b???????????1????????????????????} with (``iff_exp``); \
    wildcard bins BIT21_1 = {32'b??????????1?????????????????????} with (``iff_exp``); \
    wildcard bins BIT22_1 = {32'b?????????1??????????????????????} with (``iff_exp``); \
    wildcard bins BIT23_1 = {32'b????????1???????????????????????} with (``iff_exp``); \
    wildcard bins BIT24_1 = {32'b???????1????????????????????????} with (``iff_exp``); \
    wildcard bins BIT25_1 = {32'b??????1?????????????????????????} with (``iff_exp``); \
    wildcard bins BIT26_1 = {32'b?????1??????????????????????????} with (``iff_exp``); \
    wildcard bins BIT27_1 = {32'b????1???????????????????????????} with (``iff_exp``); \
    wildcard bins BIT28_1 = {32'b???1????????????????????????????} with (``iff_exp``); \
    wildcard bins BIT29_1 = {32'b??1?????????????????????????????} with (``iff_exp``); \
    wildcard bins BIT30_1 = {32'b?1??????????????????????????????} with (``iff_exp``); \
    wildcard bins BIT31_1 = {32'b1???????????????????????????????} with (``iff_exp``); \
}

`define CVXIF_CP_BITWISE(name, field, iff_exp) \
``name``: coverpoint(``field``) iff (``iff_exp``) { \
    wildcard bins BIT0_0  = {32'b???????????????????????????????0}; \
    wildcard bins BIT1_0  = {32'b??????????????????????????????0?}; \
    wildcard bins BIT2_0  = {32'b?????????????????????????????0??}; \
    wildcard bins BIT3_0  = {32'b????????????????????????????0???}; \
    wildcard bins BIT4_0  = {32'b???????????????????????????0????}; \
    wildcard bins BIT5_0  = {32'b??????????????????????????0?????}; \
    wildcard bins BIT6_0  = {32'b?????????????????????????0??????}; \
    wildcard bins BIT7_0  = {32'b????????????????????????0???????}; \
    wildcard bins BIT8_0  = {32'b???????????????????????0????????}; \
    wildcard bins BIT9_0  = {32'b??????????????????????0?????????}; \
    wildcard bins BIT10_0 = {32'b?????????????????????0??????????}; \
    wildcard bins BIT11_0 = {32'b????????????????????0???????????}; \
    wildcard bins BIT12_0 = {32'b???????????????????0????????????}; \
    wildcard bins BIT13_0 = {32'b??????????????????0?????????????}; \
    wildcard bins BIT14_0 = {32'b?????????????????0??????????????}; \
    wildcard bins BIT15_0 = {32'b????????????????0???????????????}; \
    wildcard bins BIT16_0 = {32'b???????????????0????????????????}; \
    wildcard bins BIT17_0 = {32'b??????????????0?????????????????}; \
    wildcard bins BIT18_0 = {32'b?????????????0??????????????????}; \
    wildcard bins BIT19_0 = {32'b????????????0???????????????????}; \
    wildcard bins BIT20_0 = {32'b???????????0????????????????????}; \
    wildcard bins BIT21_0 = {32'b??????????0?????????????????????}; \
    wildcard bins BIT22_0 = {32'b?????????0??????????????????????}; \
    wildcard bins BIT23_0 = {32'b????????0???????????????????????}; \
    wildcard bins BIT24_0 = {32'b???????0????????????????????????}; \
    wildcard bins BIT25_0 = {32'b??????0?????????????????????????}; \
    wildcard bins BIT26_0 = {32'b?????0??????????????????????????}; \
    wildcard bins BIT27_0 = {32'b????0???????????????????????????}; \
    wildcard bins BIT28_0 = {32'b???0????????????????????????????}; \
    wildcard bins BIT29_0 = {32'b??0?????????????????????????????}; \
    wildcard bins BIT30_0 = {32'b?0??????????????????????????????}; \
    wildcard bins BIT31_0 = {32'b0???????????????????????????????}; \
    wildcard bins BIT0_1  = {32'b???????????????????????????????1}; \
    wildcard bins BIT1_1  = {32'b??????????????????????????????1?}; \
    wildcard bins BIT2_1  = {32'b?????????????????????????????1??}; \
    wildcard bins BIT3_1  = {32'b????????????????????????????1???}; \
    wildcard bins BIT4_1  = {32'b???????????????????????????1????}; \
    wildcard bins BIT5_1  = {32'b??????????????????????????1?????}; \
    wildcard bins BIT6_1  = {32'b?????????????????????????1??????}; \
    wildcard bins BIT7_1  = {32'b????????????????????????1???????}; \
    wildcard bins BIT8_1  = {32'b???????????????????????1????????}; \
    wildcard bins BIT9_1  = {32'b??????????????????????1?????????}; \
    wildcard bins BIT10_1 = {32'b?????????????????????1??????????}; \
    wildcard bins BIT11_1 = {32'b????????????????????1???????????}; \
    wildcard bins BIT12_1 = {32'b???????????????????1????????????}; \
    wildcard bins BIT13_1 = {32'b??????????????????1?????????????}; \
    wildcard bins BIT14_1 = {32'b?????????????????1??????????????}; \
    wildcard bins BIT15_1 = {32'b????????????????1???????????????}; \
    wildcard bins BIT16_1 = {32'b???????????????1????????????????}; \
    wildcard bins BIT17_1 = {32'b??????????????1?????????????????}; \
    wildcard bins BIT18_1 = {32'b?????????????1??????????????????}; \
    wildcard bins BIT19_1 = {32'b????????????1???????????????????}; \
    wildcard bins BIT20_1 = {32'b???????????1????????????????????}; \
    wildcard bins BIT21_1 = {32'b??????????1?????????????????????}; \
    wildcard bins BIT22_1 = {32'b?????????1??????????????????????}; \
    wildcard bins BIT23_1 = {32'b????????1???????????????????????}; \
    wildcard bins BIT24_1 = {32'b???????1????????????????????????}; \
    wildcard bins BIT25_1 = {32'b??????1?????????????????????????}; \
    wildcard bins BIT26_1 = {32'b?????1??????????????????????????}; \
    wildcard bins BIT27_1 = {32'b????1???????????????????????????}; \
    wildcard bins BIT28_1 = {32'b???1????????????????????????????}; \
    wildcard bins BIT29_1 = {32'b??1?????????????????????????????}; \
    wildcard bins BIT30_1 = {32'b?1??????????????????????????????}; \
    wildcard bins BIT31_1 = {32'b1???????????????????????????????}; \
}

`endif // __UVMA_CVXIF_MACROS_SV__
