// ----------------------------------------------------------------------------
//Copyright 2023 CEA*
//*Commissariat a l'Energie Atomique et aux Energies Alternatives (CEA)
//
//Licensed under the Apache License, Version 2.0 (the "License");
//you may not use this file except in compliance with the License.
//You may obtain a copy of the License at
//
//    http://www.apache.org/licenses/LICENSE-2.0
//
//Unless required by applicable law or agreed to in writing, software
//distributed under the License is distributed on an "AS IS" BASIS,
//WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//See the License for the specific language governing permissions and
//limitations under the License.
//[END OF HEADER]
// ----------------------------------------------------------------------------
//  Description :
//
//
// ----------------------------------------------------------------------------

package test_pkg;

    import uvm_pkg::*;
    import uvma_axi_pkg::*;
    import dut_env_pkg::*;
    `include "uvm_macros.svh";
    `include "base_test_c.svh";
    `include "bursty_test_c.svh";


endpackage : test_pkg


