// Copyright 2022 Thales DIS SAS
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
// You may obtain a copy of the License at https://solderpad.org/licenses/
//
// Original Author: Alae Eddine EZ ZEJJARI (alae-eddine.ez-zejjari@external.thalesgroup.com)
// Co-Author: Abdelaali Khardazi

/**** AXI4 slave sequencer  ****/

`ifndef __UVMA_AXI_B_SQR_SV__
`define __UVMA_AXI_B_SQR_SV__

class uvma_axi_b_sqr_c extends uvm_sequencer#(uvma_axi_b_item_c);

   `uvm_component_utils(uvma_axi_b_sqr_c)

   uvm_analysis_export   #(uvma_axi_b_item_c)    b_resp_export;
   uvm_tlm_analysis_fifo #(uvma_axi_b_item_c)    b_resp_fifo;

   function new(string name = "uvma_axi_b_sqr_c", uvm_component parent = null);
      super.new(name, parent);
      this.b_resp_export = new("b_resp_export", this);
      this.b_resp_fifo   = new("b_resp_fifo", this);
   endfunction

   function void build_phase(uvm_phase phase);
      super.build_phase(phase);
   endfunction

   function void connect_phase(uvm_phase phase);
      super.connect_phase(phase);
      this.b_resp_export.connect(this.b_resp_fifo.analysis_export);       // Connect analysis export direct to fifo B channels
   endfunction

endclass

`endif
