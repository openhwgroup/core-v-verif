//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
// 
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


    c_sext_b_cg = new(); c_sext_b_cg.set_inst_name("obj_c_sext_b");
    c_zext_h_cg = new(); c_zext_h_cg.set_inst_name("obj_c_zext_h");
    c_sext_h_cg = new(); c_sext_h_cg.set_inst_name("obj_c_sext_h");


