// XPULP Instructions here:
    CV_LB,
    CV_LH,
    CV_LW,
    CV_ELW,
    CV_LBU,
    CV_LHU,
    CV_SB,
    CV_SH,
    CV_SW,
    CV_START,
    CV_STARTI,
    CV_END,
    CV_ENDI,
    CV_COUNT,
    CV_COUNTI,
    CV_SETUP,
    CV_SETUPI,
    CV_BEQIMM,
    CV_BNEIMM,
    CV_EXTRACT,
    CV_EXTRACTU,
    CV_EXTRACTR,
    CV_EXTRACTUR,
    CV_INSERT,
    CV_INSERTR,
    CV_BCLR,
    CV_BCLRR,
    CV_BSET,
    CV_BSETR,
    CV_BITREV,
    CV_ROR,
    CV_FF1,
    CV_FL1,
    CV_CLB,
    CV_CNT,
    CV_ABS,
    CV_SLE,
    CV_SLEU,
    CV_MIN,
    CV_MINU,
    CV_MAX,
    CV_MAXU,
    CV_EXTHS,
    CV_EXTHZ,
    CV_EXTBS,
    CV_EXTBZ,
    CV_CLIP,
    CV_CLIPU,
    CV_CLIPR,
    CV_CLIPUR,
    CV_ADDNR,
    CV_ADDUNR,
    CV_ADDRNR,
    CV_ADDURNR,
    CV_SUBNR,
    CV_SUBUNR,
    CV_SUBRNR,
    CV_SUBURNR,
    CV_ADDN,
    CV_ADDUN,
    CV_ADDRN,
    CV_ADDURN,
    CV_SUBN,
    CV_SUBUN,
    CV_SUBRN,
    CV_SUBURN,
    CV_MAC,
    CV_MSU,
    CV_MULSN,
    CV_MULHHSN,
    CV_MULSRN,
    CV_MULHHSRN,
    CV_MULUN,
    CV_MULHHUN,
    CV_MULURN,
    CV_MULHHURN,
    CV_MACSN,
    CV_MACHHSN,
    CV_MACSRN,
    CV_MACHHSRN,
    CV_MACUN,
    CV_MACHHUN,
    CV_MACURN,
    CV_MACHHURN,
    CV_ADD_H,
    CV_ADD_B,
    CV_ADD_SC_H,
    CV_ADD_SC_B,
    CV_ADD_SCI_H,
    CV_ADD_SCI_B,
    CV_SUB_H,
    CV_SUB_B,
    CV_SUB_SC_H,
    CV_SUB_SC_B,
    CV_SUB_SCI_H,
    CV_SUB_SCI_B,
    CV_AVG_H,
    CV_AVG_B,
    CV_AVG_SC_H,
    CV_AVG_SC_B,
    CV_AVG_SCI_H,
    CV_AVG_SCI_B,
    CV_AVGU_H,
    CV_AVGU_B,
    CV_AVGU_SC_H,
    CV_AVGU_SC_B,
    CV_AVGU_SCI_H,
    CV_AVGU_SCI_B,
    CV_MIN_H,
    CV_MIN_B,
    CV_MIN_SC_H,
    CV_MIN_SC_B,
    CV_MIN_SCI_H,
    CV_MIN_SCI_B,
    CV_MINU_H,
    CV_MINU_B,
    CV_MINU_SC_H,
    CV_MINU_SC_B,
    CV_MINU_SCI_H,
    CV_MINU_SCI_B,
    CV_MAX_H,
    CV_MAX_B,
    CV_MAX_SC_H,
    CV_MAX_SC_B,
    CV_MAX_SCI_H,
    CV_MAX_SCI_B,
    CV_MAXU_H,
    CV_MAXU_B,
    CV_MAXU_SC_H,
    CV_MAXU_SC_B,
    CV_MAXU_SCI_H,
    CV_MAXU_SCI_B,
    CV_SRL_H,
    CV_SRL_B,
    CV_SRL_SC_H,
    CV_SRL_SC_B,
    CV_SRL_SCI_H,
    CV_SRL_SCI_B,
    CV_SRA_H,
    CV_SRA_B,
    CV_SRA_SC_H,
    CV_SRA_SC_B,
    CV_SRA_SCI_H,
    CV_SRA_SCI_B,
    CV_SLL_H,
    CV_SLL_B,
    CV_SLL_SC_H,
    CV_SLL_SC_B,
    CV_SLL_SCI_H,
    CV_SLL_SCI_B,
    CV_OR_H,
    CV_OR_B,
    CV_OR_SC_H,
    CV_OR_SC_B,
    CV_OR_SCI_H,
    CV_OR_SCI_B,
    CV_XOR_H,
    CV_XOR_B,
    CV_XOR_SC_H,
    CV_XOR_SC_B,
    CV_XOR_SCI_H,
    CV_XOR_SCI_B,
    CV_AND_H,
    CV_AND_B,
    CV_AND_SC_H,
    CV_AND_SC_B,
    CV_AND_SCI_H,
    CV_AND_SCI_B,
    CV_ABS_H,
    CV_ABS_B,
    CV_DOTUP_H,
    CV_DOTUP_B,
    CV_DOTUP_SC_H,
    CV_DOTUP_SC_B,
    CV_DOTUP_SCI_H,
    CV_DOTUP_SCI_B,
    CV_DOTUSP_H,
    CV_DOTUSP_B,
    CV_DOTUSP_SC_H,
    CV_DOTUSP_SC_B,
    CV_DOTUSP_SCI_H,
    CV_DOTUSP_SCI_B,
    CV_DOTSP_H,
    CV_DOTSP_B,
    CV_DOTSP_SC_H,
    CV_DOTSP_SC_B,
    CV_DOTSP_SCI_H,
    CV_DOTSP_SCI_B,
    CV_SDOTUP_H,
    CV_SDOTUP_B,
    CV_SDOTUP_SC_H,
    CV_SDOTUP_SC_B,
    CV_SDOTUP_SCI_H,
    CV_SDOTUP_SCI_B,
    CV_SDOTUSP_H,
    CV_SDOTUSP_B,
    CV_SDOTUSP_SC_H,
    CV_SDOTUSP_SC_B,
    CV_SDOTUSP_SCI_H,
    CV_SDOTUSP_SCI_B,
    CV_SDOTSP_H,
    CV_SDOTSP_B,
    CV_SDOTSP_SC_H,
    CV_SDOTSP_SC_B,
    CV_SDOTSP_SCI_H,
    CV_SDOTSP_SCI_B,
    CV_EXTRACT_H,
    CV_EXTRACT_B,
    CV_EXTRACTU_H,
    CV_EXTRACTU_B,
    CV_INSERT_H,
    CV_INSERT_B,
    CV_SHUFFLE_H,
    CV_SHUFFLE_B,
    CV_SHUFFLE_SCI_H,
    CV_SHUFFLEI0_SCI_B,
    CV_SHUFFLEI1_SCI_B,
    CV_SHUFFLEI2_SCI_B,
    CV_SHUFFLEI3_SCI_B,
    CV_SHUFFLE2_H,
    CV_SHUFFLE2_B,
    CV_PACK,
    CV_PACK_H,
    CV_PACKHI_B,
    CV_PACKLO_B,
    CV_CMPEQ_H,
    CV_CMPEQ_B,
    CV_CMPEQ_SC_H,
    CV_CMPEQ_SC_B,
    CV_CMPEQ_SCI_H,
    CV_CMPEQ_SCI_B,
    CV_CMPNE_H,
    CV_CMPNE_B,
    CV_CMPNE_SC_H,
    CV_CMPNE_SC_B,
    CV_CMPNE_SCI_H,
    CV_CMPNE_SCI_B,
    CV_CMPGT_H,
    CV_CMPGT_B,
    CV_CMPGT_SC_H,
    CV_CMPGT_SC_B,
    CV_CMPGT_SCI_H,
    CV_CMPGT_SCI_B,
    CV_CMPGE_H,
    CV_CMPGE_B,
    CV_CMPGE_SC_H,
    CV_CMPGE_SC_B,
    CV_CMPGE_SCI_H,
    CV_CMPGE_SCI_B,
    CV_CMPLT_H,
    CV_CMPLT_B,
    CV_CMPLT_SC_H,
    CV_CMPLT_SC_B,
    CV_CMPLT_SCI_H,
    CV_CMPLT_SCI_B,
    CV_CMPLE_H,
    CV_CMPLE_B,
    CV_CMPLE_SC_H,
    CV_CMPLE_SC_B,
    CV_CMPLE_SCI_H,
    CV_CMPLE_SCI_B,
    CV_CMPGTU_H,
    CV_CMPGTU_B,
    CV_CMPGTU_SC_H,
    CV_CMPGTU_SC_B,
    CV_CMPGTU_SCI_H,
    CV_CMPGTU_SCI_B,
    CV_CMPGEU_H,
    CV_CMPGEU_B,
    CV_CMPGEU_SC_H,
    CV_CMPGEU_SC_B,
    CV_CMPGEU_SCI_H,
    CV_CMPGEU_SCI_B,
    CV_CMPLTU_H,
    CV_CMPLTU_B,
    CV_CMPLTU_SC_H,
    CV_CMPLTU_SC_B,
    CV_CMPLTU_SCI_H,
    CV_CMPLTU_SCI_B,
    CV_CMPLEU_H,
    CV_CMPLEU_B,
    CV_CMPLEU_SC_H,
    CV_CMPLEU_SC_B,
    CV_CMPLEU_SCI_H,
    CV_CMPLEU_SCI_B,
    CV_CPLXMUL_R,
    CV_CPLXMUL_I,
    CV_CPLXMUL_R_DIV2,
    CV_CPLXMUL_I_DIV2,
    CV_CPLXMUL_R_DIV4,
    CV_CPLXMUL_I_DIV4,
    CV_CPLXMUL_R_DIV8,
    CV_CPLXMUL_I_DIV8,
    CV_CPLXCONJ,
    CV_SUBROTMJ,
    CV_SUBROTMJ_DIV2,
    CV_SUBROTMJ_DIV4,
    CV_SUBROTMJ_DIV8,
    CV_ADD_DIV2,
    CV_ADD_DIV4,
    CV_ADD_DIV8,
    CV_SUB_DIV2,
    CV_SUB_DIV4,
    CV_SUB_DIV8,
