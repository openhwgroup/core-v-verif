//
// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2020 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//


`ifndef __UVMT_CV32E40S_TB_SV__
`define __UVMT_CV32E40S_TB_SV__

/**
 * Module encapsulating the CV32E40S DUT wrapper, and associated SV interfaces.
 * Also provide UVM environment entry and exit points.
 */
`default_nettype none
module uvmt_cv32e40s_tb;

   import uvm_pkg::*;
   import cv32e40s_pkg::*;
   import uvmt_cv32e40s_base_test_pkg::*;
   import uvmt_cv32e40s_pkg::*;
   `ifndef FORMAL
   import rvviApiPkg::*;
   `endif

   // Capture regs for test status from Virtual Peripheral in dut_wrap.mem_i
   bit        tp;
   bit        tf;
   bit        evalid;
   bit [31:0] evalue;

   // Agent interfaces
   uvma_clknrst_if_t            clknrst_if(); // clock and resets from the clknrst agent
   uvma_clknrst_if_t            clknrst_if_iss();
   uvma_debug_if_t              debug_if();
   uvma_wfe_wu_if_t             wfe_wu_if();
   uvma_interrupt_if_t          interrupt_if();
   uvma_clic_if_t#(
     .CLIC_ID_WIDTH(uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC_ID_WIDTH)
   ) clic_if();
   uvma_obi_memory_if_t #(
     .ADDR_WIDTH  (ENV_PARAM_INSTR_ADDR_WIDTH),
     .DATA_WIDTH  (ENV_PARAM_INSTR_DATA_WIDTH),
     .ACHK_WIDTH  (ENV_PARAM_INSTR_ACHK_WIDTH),
     .RCHK_WIDTH  (ENV_PARAM_INSTR_RCHK_WIDTH)
   ) obi_instr_if (
     .clk     (clknrst_if.clk),
     .reset_n (clknrst_if.reset_n)
   );

   uvma_obi_memory_if_t #(
     .ADDR_WIDTH  (ENV_PARAM_DATA_ADDR_WIDTH),
     .DATA_WIDTH  (ENV_PARAM_DATA_DATA_WIDTH),
     .ACHK_WIDTH  (ENV_PARAM_DATA_ACHK_WIDTH),
     .RCHK_WIDTH  (ENV_PARAM_DATA_RCHK_WIDTH)
   ) obi_data_if(
     .clk(clknrst_if.clk),
     .reset_n(clknrst_if.reset_n)
   );
   uvma_fencei_if_t               fencei_if(
     .clk(clknrst_if.clk),
     .reset_n(clknrst_if.reset_n)
   );

   // DUT Wrapper Interfaces
   uvmt_cv32e40s_vp_status_if_t     vp_status_if(.tests_passed(),
                                                 .tests_failed(),
                                                 .exit_valid(),
                                                 .exit_value()); // Status information generated by the Virtual Peripherals in the DUT WRAPPER memory.
   uvme_cv32e40s_core_cntrl_if_t      core_cntrl_if();

   // RVVI SystemVerilog Interface
   `ifndef FORMAL
      rvviTrace #( .NHART(1), .RETIRE(1)) rvvi_if();
      //uvmt_imperas_dv_if_t imperas_dv_if();
      uvmt_reference_model_if_t reference_model_if();
   `endif


  // "dut_wrap"

  uvmt_cv32e40s_dut_wrap  #(
    .INSTR_ADDR_WIDTH  (ENV_PARAM_INSTR_ADDR_WIDTH),
    .INSTR_RDATA_WIDTH (ENV_PARAM_INSTR_DATA_WIDTH),
    .RAM_ADDR_WIDTH    (ENV_PARAM_RAM_ADDR_WIDTH)
  ) dut_wrap (
    .clknrst_if     (clknrst_if),
    .interrupt_if   (interrupt_if),
    .vp_status_if   (vp_status_if),
    .core_cntrl_if  (core_cntrl_if),
    .obi_instr_if   (obi_instr_if),
    .obi_data_if    (obi_data_if),
    .fencei_if      (fencei_if),
    .clic_if        (clic_if),
    .*
  );

  assign debug_if.clk     = clknrst_if.clk;
  assign debug_if.reset_n = clknrst_if.reset_n;

  // OBI Instruction agent v1.2 signal tie-offs
  assign obi_instr_if.we        = 'b0;
  assign obi_instr_if.be        = 'hf; // Always assumes 32-bit full bus reads on instruction OBI
  assign obi_instr_if.auser     = 'b0;
  assign obi_instr_if.wuser     = 'b0;
  assign obi_instr_if.aid       = 'b0;
  assign obi_instr_if.wdata     = 'b0;
  assign obi_instr_if.rready    = 1'b1;
  assign obi_instr_if.rreadypar = 1'b0;

  // OBI Data agent v1.2 signal tie-offs
  assign obi_data_if.auser     = 'b0;
  assign obi_data_if.wuser     = 'b0;
  assign obi_data_if.aid       = 'b0;
  assign obi_data_if.rready    = 1'b1;
  assign obi_data_if.rreadypar = 1'b0;

  // Connect to uvma_interrupt_if
  assign interrupt_if.clk     = clknrst_if.clk;
  assign interrupt_if.reset_n = clknrst_if.reset_n;
  assign interrupt_if.irq_id  = $bits(interrupt_if.irq_id)'(dut_wrap.cv32e40s_wrapper_i.core_i.irq_id); // cast to avoid the warning with clic (TODO: tieoff with clic instead?)
  assign interrupt_if.irq_ack = dut_wrap.cv32e40s_wrapper_i.core_i.irq_ack;

  assign clic_if.clk     = clknrst_if.clk;
  assign clic_if.reset_n = clknrst_if.reset_n;
  assign clic_if.irq_ack = dut_wrap.cv32e40s_wrapper_i.core_i.irq_ack;

  assign wfe_wu_if.clk     = clknrst_if.clk;
  assign wfe_wu_if.reset_n = clknrst_if.reset_n;

  // Connect to core_cntrl_if
  assign core_cntrl_if.b_ext = uvmt_cv32e40s_base_test_pkg::CORE_PARAM_B_EXT;
  `ifndef FORMAL
    initial begin
      core_cntrl_if.pma_cfg = new[CORE_PARAM_PMA_NUM_REGIONS];
      foreach (core_cntrl_if.pma_cfg[i]) begin
        core_cntrl_if.pma_cfg[i].word_addr_low  = CORE_PARAM_PMA_CFG[i].word_addr_low;
        core_cntrl_if.pma_cfg[i].word_addr_high = CORE_PARAM_PMA_CFG[i].word_addr_high;
        core_cntrl_if.pma_cfg[i].main           = CORE_PARAM_PMA_CFG[i].main;
        core_cntrl_if.pma_cfg[i].bufferable     = CORE_PARAM_PMA_CFG[i].bufferable;
        core_cntrl_if.pma_cfg[i].cacheable      = CORE_PARAM_PMA_CFG[i].cacheable;
        core_cntrl_if.pma_cfg[i].integrity      = CORE_PARAM_PMA_CFG[i].integrity;
      end
    end
  `endif


  // "rvfi_instr_if"

  bind cv32e40s_wrapper
    uvma_rvfi_instr_if_t#(
      uvmt_cv32e40s_base_test_pkg::ILEN,
      uvmt_cv32e40s_base_test_pkg::XLEN
    ) rvfi_instr_if(
      .clk (clk_i),
      .reset_n (rst_ni),

      .rvfi_valid (rvfi_i.rvfi_valid[0]),
      .rvfi_order (rvfi_i.rvfi_order[uvma_rvfi_pkg::ORDER_WL*0+:uvma_rvfi_pkg::ORDER_WL]),
      .rvfi_insn (rvfi_i.rvfi_insn[uvmt_cv32e40s_base_test_pkg::ILEN*0+:uvmt_cv32e40s_base_test_pkg::ILEN]),
      .rvfi_trap (rvfi_i.rvfi_trap),
      .rvfi_halt (rvfi_i.rvfi_halt[0]),
      .rvfi_intr (rvfi_i.rvfi_intr),
      .rvfi_dbg (rvfi_i.rvfi_dbg),
      .rvfi_dbg_mode (rvfi_i.rvfi_dbg_mode),
      .rvfi_nmip (rvfi_i.rvfi_nmip),
      .rvfi_mode (rvfi_i.rvfi_mode[uvma_rvfi_pkg::MODE_WL*0+:uvma_rvfi_pkg::MODE_WL]),
      .rvfi_ixl (rvfi_i.rvfi_ixl[uvma_rvfi_pkg::IXL_WL*0+:uvma_rvfi_pkg::IXL_WL]),
      .rvfi_pc_rdata (rvfi_i.rvfi_pc_rdata[uvmt_cv32e40s_base_test_pkg::XLEN*0+:uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_pc_wdata (rvfi_i.rvfi_pc_wdata[uvmt_cv32e40s_base_test_pkg::XLEN*0+:uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_rs1_addr (rvfi_i.rvfi_rs1_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
      .rvfi_rs1_rdata (rvfi_i.rvfi_rs1_rdata[uvmt_cv32e40s_base_test_pkg::XLEN*0+:uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_rs2_addr (rvfi_i.rvfi_rs2_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
      .rvfi_rs2_rdata (rvfi_i.rvfi_rs2_rdata[uvmt_cv32e40s_base_test_pkg::XLEN*0+:uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_rs3_addr ('0),
      .rvfi_rs3_rdata ('0),
      .rvfi_rd1_addr (rvfi_i.rvfi_rd_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
      .rvfi_rd1_wdata (rvfi_i.rvfi_rd_wdata[uvmt_cv32e40s_base_test_pkg::XLEN*0+:uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_rd2_addr ('0),
      .rvfi_rd2_wdata ('0),
      .rvfi_gpr_rdata (rvfi_i.rvfi_gpr_rdata[32*uvmt_cv32e40s_base_test_pkg::XLEN*0  +:32*uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_gpr_rmask (rvfi_i.rvfi_gpr_rmask[32*0  +:32]),
      .rvfi_gpr_wdata (rvfi_i.rvfi_gpr_wdata[32*uvmt_cv32e40s_base_test_pkg::XLEN*0  +:32*uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_gpr_wmask (rvfi_i.rvfi_gpr_wmask[32*0  +:32]),
      .rvfi_mem_addr (rvfi_i.rvfi_mem_addr[  uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_mem_rdata (rvfi_i.rvfi_mem_rdata[uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_mem_rmask (rvfi_i.rvfi_mem_rmask[uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN/8*0  +:uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN/8]),
      .rvfi_mem_wdata (rvfi_i.rvfi_mem_wdata[uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN]),
      .rvfi_mem_wmask (rvfi_i.rvfi_mem_wmask[uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN/8*0  +:uvma_rvfi_pkg::NMEM*uvmt_cv32e40s_base_test_pkg::XLEN/8]),
      .rvfi_instr_prot (rvfi_i.rvfi_instr_prot),
      .rvfi_instr_memtype (rvfi_i.rvfi_instr_memtype),
      .rvfi_instr_dbg (rvfi_i.rvfi_instr_dbg),
      .rvfi_mem_prot (rvfi_i.rvfi_mem_prot),
      .rvfi_mem_exokay (rvfi_i.rvfi_mem_exokay),
      .rvfi_mem_err (rvfi_i.rvfi_mem_err),
      .rvfi_mem_atop (rvfi_i.rvfi_mem_atop),
      .rvfi_mem_memtype (rvfi_i.rvfi_mem_memtype),
      .rvfi_mem_dbg (rvfi_i.rvfi_mem_dbg)
    );

  // RVFI CSR binds
  `RVFI_CSR_BIND(cpuctrl)
  `RVFI_CSR_BIND(jvt)
  `RVFI_CSR_BIND(marchid)
  `RVFI_CSR_BIND(mcause)
  `RVFI_CSR_BIND(mcounteren)
  `RVFI_CSR_BIND(mcountinhibit)
  `RVFI_CSR_BIND(mcycle)
  `RVFI_CSR_BIND(mcycleh)
  `RVFI_CSR_BIND(menvcfg)
  `RVFI_CSR_BIND(menvcfgh)
  `RVFI_CSR_BIND(mepc)
  `RVFI_CSR_BIND(mhartid)
  `RVFI_CSR_BIND(mie)
  `RVFI_CSR_BIND(mimpid)
  `RVFI_CSR_BIND(minstret)
  `RVFI_CSR_BIND(minstreth)
  `RVFI_CSR_BIND(mip)
  `RVFI_CSR_BIND(misa)
  `RVFI_CSR_BIND(mscratch)
  `RVFI_CSR_BIND(mstateen0)
  `RVFI_CSR_BIND(mstateen1)
  `RVFI_CSR_BIND(mstateen2)
  `RVFI_CSR_BIND(mstateen3)
  `RVFI_CSR_BIND(mstateen0h)
  `RVFI_CSR_BIND(mstateen1h)
  `RVFI_CSR_BIND(mstateen2h)
  `RVFI_CSR_BIND(mstateen3h)
  `RVFI_CSR_BIND(mstatus)
  `RVFI_CSR_BIND(mstatush)
  `RVFI_CSR_BIND(mtval)
  `RVFI_CSR_BIND(mtvec)
  `RVFI_CSR_BIND(mvendorid)
  `RVFI_CSR_BIND(mseccfg)
  `RVFI_CSR_BIND(mseccfgh)

  `RVFI_CSR_BIND(dcsr)
  `RVFI_CSR_BIND(dpc)
  `RVFI_CSR_BIND(tselect)
  `RVFI_CSR_BIND(tinfo)

  `RVFI_CSR_IDX_BIND(mhpmcounter,,3)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,4)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,5)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,6)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,7)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,8)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,9)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,10)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,11)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,12)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,13)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,14)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,15)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,16)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,17)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,18)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,19)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,20)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,21)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,22)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,23)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,24)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,25)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,26)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,27)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,28)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,29)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,30)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,31)

  `RVFI_CSR_IDX_BIND(pmpcfg,,0)
  `RVFI_CSR_IDX_BIND(pmpcfg,,1)
  `RVFI_CSR_IDX_BIND(pmpcfg,,2)
  `RVFI_CSR_IDX_BIND(pmpcfg,,3)
  `RVFI_CSR_IDX_BIND(pmpcfg,,4)
  `RVFI_CSR_IDX_BIND(pmpcfg,,5)
  `RVFI_CSR_IDX_BIND(pmpcfg,,6)
  `RVFI_CSR_IDX_BIND(pmpcfg,,7)
  `RVFI_CSR_IDX_BIND(pmpcfg,,8)
  `RVFI_CSR_IDX_BIND(pmpcfg,,9)
  `RVFI_CSR_IDX_BIND(pmpcfg,,10)
  `RVFI_CSR_IDX_BIND(pmpcfg,,11)
  `RVFI_CSR_IDX_BIND(pmpcfg,,12)
  `RVFI_CSR_IDX_BIND(pmpcfg,,13)
  `RVFI_CSR_IDX_BIND(pmpcfg,,14)
  `RVFI_CSR_IDX_BIND(pmpcfg,,15)

  `RVFI_CSR_IDX_BIND(pmpaddr,,0)
  `RVFI_CSR_IDX_BIND(pmpaddr,,1)
  `RVFI_CSR_IDX_BIND(pmpaddr,,2)
  `RVFI_CSR_IDX_BIND(pmpaddr,,3)
  `RVFI_CSR_IDX_BIND(pmpaddr,,4)
  `RVFI_CSR_IDX_BIND(pmpaddr,,5)
  `RVFI_CSR_IDX_BIND(pmpaddr,,6)
  `RVFI_CSR_IDX_BIND(pmpaddr,,7)
  `RVFI_CSR_IDX_BIND(pmpaddr,,8)
  `RVFI_CSR_IDX_BIND(pmpaddr,,9)
  `RVFI_CSR_IDX_BIND(pmpaddr,,10)
  `RVFI_CSR_IDX_BIND(pmpaddr,,11)
  `RVFI_CSR_IDX_BIND(pmpaddr,,12)
  `RVFI_CSR_IDX_BIND(pmpaddr,,13)
  `RVFI_CSR_IDX_BIND(pmpaddr,,14)
  `RVFI_CSR_IDX_BIND(pmpaddr,,15)
  `RVFI_CSR_IDX_BIND(pmpaddr,,16)
  `RVFI_CSR_IDX_BIND(pmpaddr,,17)
  `RVFI_CSR_IDX_BIND(pmpaddr,,18)
  `RVFI_CSR_IDX_BIND(pmpaddr,,19)
  `RVFI_CSR_IDX_BIND(pmpaddr,,20)
  `RVFI_CSR_IDX_BIND(pmpaddr,,21)
  `RVFI_CSR_IDX_BIND(pmpaddr,,22)
  `RVFI_CSR_IDX_BIND(pmpaddr,,23)
  `RVFI_CSR_IDX_BIND(pmpaddr,,24)
  `RVFI_CSR_IDX_BIND(pmpaddr,,25)
  `RVFI_CSR_IDX_BIND(pmpaddr,,26)
  `RVFI_CSR_IDX_BIND(pmpaddr,,27)
  `RVFI_CSR_IDX_BIND(pmpaddr,,28)
  `RVFI_CSR_IDX_BIND(pmpaddr,,29)
  `RVFI_CSR_IDX_BIND(pmpaddr,,30)
  `RVFI_CSR_IDX_BIND(pmpaddr,,31)
  `RVFI_CSR_IDX_BIND(pmpaddr,,32)
  `RVFI_CSR_IDX_BIND(pmpaddr,,33)
  `RVFI_CSR_IDX_BIND(pmpaddr,,34)
  `RVFI_CSR_IDX_BIND(pmpaddr,,35)
  `RVFI_CSR_IDX_BIND(pmpaddr,,36)
  `RVFI_CSR_IDX_BIND(pmpaddr,,37)
  `RVFI_CSR_IDX_BIND(pmpaddr,,38)
  `RVFI_CSR_IDX_BIND(pmpaddr,,39)
  `RVFI_CSR_IDX_BIND(pmpaddr,,40)
  `RVFI_CSR_IDX_BIND(pmpaddr,,41)
  `RVFI_CSR_IDX_BIND(pmpaddr,,42)
  `RVFI_CSR_IDX_BIND(pmpaddr,,43)
  `RVFI_CSR_IDX_BIND(pmpaddr,,44)
  `RVFI_CSR_IDX_BIND(pmpaddr,,45)
  `RVFI_CSR_IDX_BIND(pmpaddr,,46)
  `RVFI_CSR_IDX_BIND(pmpaddr,,47)
  `RVFI_CSR_IDX_BIND(pmpaddr,,48)
  `RVFI_CSR_IDX_BIND(pmpaddr,,49)
  `RVFI_CSR_IDX_BIND(pmpaddr,,50)
  `RVFI_CSR_IDX_BIND(pmpaddr,,51)
  `RVFI_CSR_IDX_BIND(pmpaddr,,52)
  `RVFI_CSR_IDX_BIND(pmpaddr,,53)
  `RVFI_CSR_IDX_BIND(pmpaddr,,54)
  `RVFI_CSR_IDX_BIND(pmpaddr,,55)
  `RVFI_CSR_IDX_BIND(pmpaddr,,56)
  `RVFI_CSR_IDX_BIND(pmpaddr,,57)
  `RVFI_CSR_IDX_BIND(pmpaddr,,58)
  `RVFI_CSR_IDX_BIND(pmpaddr,,59)
  `RVFI_CSR_IDX_BIND(pmpaddr,,60)
  `RVFI_CSR_IDX_BIND(pmpaddr,,61)
  `RVFI_CSR_IDX_BIND(pmpaddr,,62)
  `RVFI_CSR_IDX_BIND(pmpaddr,,63)

  `RVFI_CSR_IDX_BIND(mhpmevent,,3)
  `RVFI_CSR_IDX_BIND(mhpmevent,,4)
  `RVFI_CSR_IDX_BIND(mhpmevent,,5)
  `RVFI_CSR_IDX_BIND(mhpmevent,,6)
  `RVFI_CSR_IDX_BIND(mhpmevent,,7)
  `RVFI_CSR_IDX_BIND(mhpmevent,,8)
  `RVFI_CSR_IDX_BIND(mhpmevent,,9)
  `RVFI_CSR_IDX_BIND(mhpmevent,,10)
  `RVFI_CSR_IDX_BIND(mhpmevent,,11)
  `RVFI_CSR_IDX_BIND(mhpmevent,,12)
  `RVFI_CSR_IDX_BIND(mhpmevent,,13)
  `RVFI_CSR_IDX_BIND(mhpmevent,,14)
  `RVFI_CSR_IDX_BIND(mhpmevent,,15)
  `RVFI_CSR_IDX_BIND(mhpmevent,,16)
  `RVFI_CSR_IDX_BIND(mhpmevent,,17)
  `RVFI_CSR_IDX_BIND(mhpmevent,,18)
  `RVFI_CSR_IDX_BIND(mhpmevent,,19)
  `RVFI_CSR_IDX_BIND(mhpmevent,,20)
  `RVFI_CSR_IDX_BIND(mhpmevent,,21)
  `RVFI_CSR_IDX_BIND(mhpmevent,,22)
  `RVFI_CSR_IDX_BIND(mhpmevent,,23)
  `RVFI_CSR_IDX_BIND(mhpmevent,,24)
  `RVFI_CSR_IDX_BIND(mhpmevent,,25)
  `RVFI_CSR_IDX_BIND(mhpmevent,,26)
  `RVFI_CSR_IDX_BIND(mhpmevent,,27)
  `RVFI_CSR_IDX_BIND(mhpmevent,,28)
  `RVFI_CSR_IDX_BIND(mhpmevent,,29)
  `RVFI_CSR_IDX_BIND(mhpmevent,,30)
  `RVFI_CSR_IDX_BIND(mhpmevent,,31)

  `RVFI_CSR_IDX_BIND(mhpmcounter,h,3)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,4)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,5)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,6)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,7)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,8)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,9)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,10)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,11)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,12)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,13)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,14)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,15)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,16)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,17)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,18)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,19)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,20)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,21)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,22)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,23)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,24)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,25)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,26)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,27)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,28)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,29)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,30)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,31)

  `RVFI_CSR_BIND(mconfigptr)
  `RVFI_CSR_BIND(secureseed0)
  `RVFI_CSR_BIND(secureseed1)
  `RVFI_CSR_BIND(secureseed2)

  if (CORE_PARAM_CLIC == 1) begin: gen_clic_rvfi_bind
    `RVFI_CSR_BIND(mintstatus)
    `RVFI_CSR_BIND(mintthresh)
    `RVFI_CSR_BIND(mnxti)
    `RVFI_CSR_BIND(mscratchcsw)
    `RVFI_CSR_BIND(mscratchcswl)
    `RVFI_CSR_BIND(mtvt)
  end : gen_clic_rvfi_bind

  // dscratch0
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if_t#(uvmt_cv32e40s_base_test_pkg::XLEN) rvfi_csr_dscratch0_if(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_dscratch_rmask[0]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_dscratch_wmask[0]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_dscratch_rdata[0]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_dscratch_wdata[0])
    );


  // dscratch1
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if_t#(uvmt_cv32e40s_base_test_pkg::XLEN) rvfi_csr_dscratch1_if(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_dscratch_rmask[1]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_dscratch_wmask[1]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_dscratch_rdata[1]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_dscratch_wdata[1])
    );

  // tdata1
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if_t#(uvmt_cv32e40s_base_test_pkg::XLEN) rvfi_csr_tdata1_if(.clk(clk_i),
                                                                  .reset_n(rst_ni),
                                                                  .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[1]),
                                                                  .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[1]),
                                                                  .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[1]),
                                                                  .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[1])
    );

  // tdata2
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if_t#(uvmt_cv32e40s_base_test_pkg::XLEN) rvfi_csr_tdata2_if(.clk(clk_i),
                                                                  .reset_n(rst_ni),
                                                                  .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[2]),
                                                                  .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[2]),
                                                                  .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[2]),
                                                                  .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[2])
    );



  // Bind in verification modules to the design

  bind uvmt_cv32e40s_dut_wrap
    uvma_obi_memory_assert_if_wrp#(
      .ADDR_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_ADDR_WIDTH),
      .DATA_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_DATA_WIDTH),
      .AUSER_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_AUSER_WIDTH),
      .WUSER_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_WUSER_WIDTH),
      .RUSER_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_RUSER_WIDTH),
      .ID_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_ID_WIDTH),
      .ACHK_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_ACHK_WIDTH),
      .RCHK_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_INSTR_RCHK_WIDTH),
      .IS_1P2(1)
    ) obi_instr_memory_assert_i(.obi(obi_instr_if));

  bind uvmt_cv32e40s_dut_wrap
    uvma_obi_memory_assert_if_wrp#(
      .ADDR_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_ADDR_WIDTH),
      .DATA_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_DATA_WIDTH),
      .AUSER_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_AUSER_WIDTH),
      .WUSER_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_WUSER_WIDTH),
      .RUSER_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_RUSER_WIDTH),
      .ID_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_ID_WIDTH),
      .ACHK_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_ACHK_WIDTH),
      .RCHK_WIDTH(uvmt_cv32e40s_base_test_pkg::ENV_PARAM_DATA_RCHK_WIDTH),
      .IS_1P2(1)
    ) obi_data_memory_assert_i(.obi(obi_data_if));


  if (CORE_PARAM_CLIC == 0) begin: gen_interrupt_assert
    `ifndef  COREV_ASSERT_OFF
      bind cv32e40s_core
        uvmt_cv32e40s_interrupt_assert  interrupt_assert_i (
          .dcsr_step    (cs_registers_i.dcsr_q.step),
          .mcause_n     ({cs_registers_i.mcause_n.irq, cs_registers_i.mcause_n.exception_code[4:0]}),
          .mie_q        (cs_registers_i.mie_q),
          .mip          (cs_registers_i.mip_rdata),
          .mstatus_mie  (cs_registers_i.mstatus_q.mie),
          .mstatus_tw   (cs_registers_i.mstatus_q.tw),
          .mtvec_mode_q (cs_registers_i.mtvec_q.mode),

          .if_stage_instr_rdata_i  (if_stage_i.m_c_obi_instr_if.resp_payload.rdata),
          .if_stage_instr_req_o    (if_stage_i.m_c_obi_instr_if.s_req.req),
          .if_stage_instr_rvalid_i (if_stage_i.m_c_obi_instr_if.s_rvalid.rvalid),
          .alignbuf_outstanding    (if_stage_i.prefetch_unit_i.alignment_buffer_i.outstanding_cnt_q),

          .ex_stage_instr_valid (ex_stage_i.id_ex_pipe_i.instr_valid),

          .wb_kill                   (ctrl_fsm.kill_wb),
          .wb_stage_instr_err_i      (wb_stage_i.ex_wb_pipe_i.instr.bus_resp.err),
          .wb_stage_instr_mpu_status (wb_stage_i.ex_wb_pipe_i.instr.mpu_status),
          .wb_stage_instr_rdata_i    (wb_stage_i.ex_wb_pipe_i.instr.bus_resp.rdata),
          .wb_stage_instr_valid_i    (wb_stage_i.ex_wb_pipe_i.instr_valid),
          .wb_trigger                (controller_i.controller_fsm_i.trigger_match_in_wb),
          .wb_valid                  (wb_stage_i.wb_valid),

          .branch_taken_ex (controller_i.controller_fsm_i.branch_taken_ex),
          .debug_mode_q    (controller_i.controller_fsm_i.debug_mode_q),
          .pending_nmi     (controller_i.controller_fsm_i.pending_nmi),

          .irq_ack_o (core_i.irq_ack),
          .irq_id_o  (core_i.irq_id),

          .mpu_instr_rvalid (if_stage_i.mpu_i.core_resp_valid_o),
          .obi_instr_if     (dut_wrap.obi_instr_if),
          .obi_data_if      (dut_wrap.obi_data_if),

          .writebufstate (load_store_unit_i.write_buffer_i.state),
          .rvfi          (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
          .support_if    (cv32e40s_wrapper.support_logic_module_o_if.slave_mp),

          .*
        );
    `endif
  end : gen_interrupt_assert

  if (CORE_PARAM_CLIC == 1) begin: gen_clic_assert
    // CLIC assertions
    `ifndef  COREV_ASSERT_OFF
      bind cv32e40s_core
        uvmt_cv32e40s_clic_interrupt_assert#(
          .CLIC (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC),
          .CLIC_ID_WIDTH (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC_ID_WIDTH)
        ) clic_assert_i(
          .support_if (cv32e40s_wrapper.support_logic_module_o_if.slave_mp),
          .rvfi_if(cv32e40s_wrapper.rvfi_instr_if),
          .csr_mepc_if(cv32e40s_wrapper.rvfi_csr_mepc_if),
          .csr_mstatus_if(cv32e40s_wrapper.rvfi_csr_mstatus_if),
          .csr_mcause_if(cv32e40s_wrapper.rvfi_csr_mcause_if),
          .csr_mintthresh_if(cv32e40s_wrapper.rvfi_csr_mintthresh_if),
          .csr_mintstatus_if(cv32e40s_wrapper.rvfi_csr_mintstatus_if),
          .csr_dcsr_if(cv32e40s_wrapper.rvfi_csr_dcsr_if),

          .dpc                 (cs_registers_i.dpc_rdata),
          .mintstatus          (cs_registers_i.mintstatus_rdata),
          .mintthresh          (cs_registers_i.mintthresh_rdata),
          .mcause              (cs_registers_i.mcause_rdata),
          .mtvec               (cs_registers_i.mtvec_rdata),
          .mtvt                (cs_registers_i.mtvt_rdata),
          .mepc                (cs_registers_i.mepc_rdata),
          .mip                 (cs_registers_i.mip_rdata),
          .mie                 (cs_registers_i.mie_rdata),
          .mnxti               (cs_registers_i.mnxti_rdata),
          .mscratch            (cs_registers_i.mscratch_rdata),
          .mscratchcsw         (cs_registers_i.mscratchcsw_rdata),
          .mscratchcswl        (cs_registers_i.mscratchcswl_rdata),
          .dcsr                (cs_registers_i.dcsr_rdata),

          //Control signals:
          .pc_set              (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.pc_set),
          .pc_mux              (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.pc_mux),

          .rvfi_mepc_wdata     (rvfi_i.rvfi_csr_mepc_wdata),
          .rvfi_mepc_wmask     (rvfi_i.rvfi_csr_mepc_wmask),
          .rvfi_mepc_rdata     (rvfi_i.rvfi_csr_mepc_rdata),
          .rvfi_mepc_rmask     (rvfi_i.rvfi_csr_mepc_rmask),
          .rvfi_dpc_rdata      (rvfi_i.rvfi_csr_dpc_rdata),
          .rvfi_dpc_rmask      (rvfi_i.rvfi_csr_dpc_rmask),
          .rvfi_mscratch_rdata (rvfi_i.rvfi_csr_mscratch_rdata),
          .rvfi_mscratch_rmask (rvfi_i.rvfi_csr_mscratch_rmask),
          .rvfi_mscratch_wdata (rvfi_i.rvfi_csr_mscratch_wdata),
          .rvfi_mscratch_wmask (rvfi_i.rvfi_csr_mscratch_wmask),
          .rvfi_mcause_wdata   (rvfi_i.rvfi_csr_mcause_wdata),
          .rvfi_mcause_wmask   (rvfi_i.rvfi_csr_mcause_wmask),

          .irq_i               (core_i.irq_i),
          .irq_ack             (core_i.irq_ack),
          .fetch_enable        (core_i.fetch_enable),
          .current_priv_mode   (core_i.priv_lvl),
          .mtvec_addr_i        (core_i.mtvec_addr_i),
          // External inputs
          .clic_if             (dut_wrap.clic_if),
          // Internal sampled   variants
          .irq_id              (core_i.irq_id[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC_ID_WIDTH-1:0]),
          .irq_level           (core_i.irq_level),
          .irq_priv            (core_i.irq_priv),
          .irq_shv             (core_i.irq_shv),

          .obi_instr_req       (core_i.instr_req_o),
          .obi_instr_gnt       (core_i.instr_gnt_i),
          .obi_instr_rvalid    (core_i.instr_rvalid_i),
          .obi_instr_addr      (core_i.instr_addr_o),
          .obi_instr_rdata     (core_i.instr_rdata_i),
          .obi_instr_rready    (1'b1),
          .obi_instr_err       (core_i.instr_err_i),

          .obi_data_addr       (core_i.data_addr_o),
          .obi_data_wdata      (core_i.data_wdata_o),
          .obi_data_we         (core_i.data_we_o),
          .obi_data_be         (core_i.data_be_o),
          .obi_data_req        (core_i.data_req_o),
          .obi_data_gnt        (core_i.data_gnt_i),
          .obi_data_rvalid     (core_i.data_rvalid_i),
          .obi_data_rready     (1'b1),
          .obi_data_err        (core_i.data_err_i),

          .debug_mode          (controller_i.controller_fsm_i.debug_mode_q),
          .debug_req           (core_i.debug_req_i),
          .debug_havereset     (core_i.debug_havereset_o),
          .debug_running       (core_i.debug_running_o),
          .debug_halt_addr     (dut_wrap.cv32e40s_wrapper_i.dm_halt_addr_i),
          .debug_exc_addr      (dut_wrap.cv32e40s_wrapper_i.dm_exception_addr_i),

          .rvfi_mode           (rvfi_i.rvfi_mode),
          .rvfi_insn           (rvfi_i.rvfi_insn),
          .rvfi_intr           (rvfi_i.rvfi_intr),
          .rvfi_rs1_rdata      (rvfi_i.rvfi_rs1_rdata),
          .rvfi_rs2_rdata      (rvfi_i.rvfi_rs2_rdata),
          .rvfi_rd_wdata       (rvfi_i.rvfi_rd_wdata),
          .rvfi_valid          (rvfi_i.rvfi_valid),
          .rvfi_pc_rdata       (rvfi_i.rvfi_pc_rdata),
          .rvfi_pc_wdata       (rvfi_i.rvfi_pc_wdata),
          .rvfi_trap           (rvfi_i.rvfi_trap),
          .rvfi_dbg_mode       (rvfi_i.rvfi_dbg_mode),
          .rvfi_dbg            (rvfi_i.rvfi_dbg),

          .wu_wfe              (dut_wrap.cv32e40s_wrapper_i.wu_wfe_i),
          .core_sleep_o        (core_i.core_sleep_o),
          .*
        );
    `endif
  end : gen_clic_assert


  // User-Mode Assertions

  `ifndef  COREV_ASSERT_OFF
    bind  cv32e40s_wrapper
      uvmt_cv32e40s_umode_assert #(
        .CLIC (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC)
      ) umode_assert_i (
        .rvfi_valid    (rvfi_i.rvfi_valid),
        .rvfi_mode     (rvfi_i.rvfi_mode),
        .rvfi_order    (rvfi_i.rvfi_order),
        .rvfi_trap     (rvfi_i.rvfi_trap),
        .rvfi_intr     (rvfi_i.rvfi_intr),
        .rvfi_insn     (rvfi_i.rvfi_insn),
        .rvfi_dbg_mode (rvfi_i.rvfi_dbg_mode),
        .rvfi_dbg      (rvfi_i.rvfi_dbg),
        .rvfi_pc_rdata (rvfi_i.rvfi_pc_rdata),
        .rvfi_if       (rvfi_instr_if),

        .rvfi_csr_dcsr_rdata       (rvfi_i.rvfi_csr_dcsr_rdata),
        .rvfi_csr_mcause_rdata     (rvfi_i.rvfi_csr_mcause_rdata),
        .rvfi_csr_mcause_wdata     (rvfi_i.rvfi_csr_mcause_wdata),
        .rvfi_csr_mcause_wmask     (rvfi_i.rvfi_csr_mcause_wmask),
        .rvfi_csr_mcounteren_rdata (rvfi_i.rvfi_csr_mcounteren_rdata),
        .rvfi_csr_mie_rdata        (rvfi_i.rvfi_csr_mie_rdata),
        .rvfi_csr_mip_rdata        (rvfi_i.rvfi_csr_mip_rdata),
        .rvfi_csr_misa_rdata       (rvfi_i.rvfi_csr_misa_rdata),
        .rvfi_csr_mscratch_rdata   (rvfi_i.rvfi_csr_mscratch_rdata),
        .rvfi_csr_mscratch_rmask   (rvfi_i.rvfi_csr_mscratch_rmask),
        .rvfi_csr_mscratch_wdata   (rvfi_i.rvfi_csr_mscratch_wdata),
        .rvfi_csr_mscratch_wmask   (rvfi_i.rvfi_csr_mscratch_wmask),
        .rvfi_csr_mstateen0_rdata  (rvfi_i.rvfi_csr_mstateen0_rdata),
        .rvfi_csr_mstatus_rdata    (rvfi_i.rvfi_csr_mstatus_rdata),
        .rvfi_csr_mstatus_wdata    (rvfi_i.rvfi_csr_mstatus_wdata),
        .rvfi_csr_mstatus_wmask    (rvfi_i.rvfi_csr_mstatus_wmask),

        .mpu_iside_valid (core_i.if_stage_i.mpu_i.core_trans_valid_i),
        .mpu_iside_addr  (core_i.if_stage_i.mpu_i.core_trans_i.addr),

        .obi_iside_prot (core_i.instr_prot_o),
        .obi_dside_prot (core_i.data_prot_o),

        .*
      );
  `endif


  // User-mode Coverage

  `ifndef  COREV_ASSERT_OFF
    bind  cv32e40s_wrapper
      uvmt_cv32e40s_umode_cov  umode_cov_i (
        .rvfi_valid     (rvfi_i.rvfi_valid),
        .rvfi_trap      (rvfi_i.rvfi_trap),
        .rvfi_intr      (rvfi_i.rvfi_intr),
        .rvfi_insn      (rvfi_i.rvfi_insn),
        .rvfi_rs1_rdata (rvfi_i.rvfi_rs1_rdata),
        .rvfi_pc_rdata  (rvfi_i.rvfi_pc_rdata),
        .rvfi_mode      (rvfi_i.rvfi_mode),
        .rvfi_rd_addr   (rvfi_i.rvfi_rd_addr),
        .rvfi_dbg_mode  (rvfi_i.rvfi_dbg_mode),
        .rvfi_order     (rvfi_i.rvfi_order),
        .rvfi_mem_rmask (rvfi_i.rvfi_mem_rmask),
        .rvfi_mem_wmask (rvfi_i.rvfi_mem_wmask),

        .rvfi_csr_mstatus_rdata (rvfi_i.rvfi_csr_mstatus_rdata),
        .rvfi_csr_mstatus_rmask (rvfi_i.rvfi_csr_mstatus_rmask),
        .rvfi_csr_dcsr_rdata    (rvfi_i.rvfi_csr_dcsr_rdata),
        .rvfi_csr_dcsr_rmask    (rvfi_i.rvfi_csr_dcsr_rmask),

        .obi_iside_req  (core_i.instr_req_o),
        .obi_iside_gnt  (core_i.instr_gnt_i),
        .obi_iside_addr (core_i.instr_addr_o),
        .obi_iside_prot (core_i.instr_prot_o),

        .*
      );
  `endif


  // Fence.i assertions

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_fencei_assert #(
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG)
      ) fencei_assert_i (
        .wb_valid           (core_i.wb_stage_i.wb_valid),
        .wb_instr_valid     (core_i.ex_wb_pipe.instr_valid),
        .wb_sys_en          (core_i.ex_wb_pipe.sys_en),
        .wb_sys_fencei_insn (core_i.ex_wb_pipe.sys_fencei_insn),
        .wb_pc              (core_i.ex_wb_pipe.pc),
        .wb_rdata           (core_i.ex_wb_pipe.instr.bus_resp.rdata),
        .wb_buffer_state    (core_i.load_store_unit_i.write_buffer_i.state),

        .rvfi_if (rvfi_instr_if),

        .*
      );
  `endif


  // RVFI Asserts & Covers

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.rvfi_i
      uvmt_cv32e40s_rvfi_assert #(
        .CLIC          (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC),
        .CLIC_ID_WIDTH (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC_ID_WIDTH)
      ) rvfi_assert_i (
        .rvfi_if          (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
        .support_if       (dut_wrap.cv32e40s_wrapper_i.support_logic_module_o_if.slave_mp),
        .writebuf_ready_o (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.ready_o),
        .writebuf_valid_i (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.valid_i),
        .*
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.rvfi_i
      uvmt_cv32e40s_rvfi_cov  rvfi_cov_i (
        .rvfi_if (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
        .*
      );
  `endif


  // Core integration assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_integration_assert  integration_assert_i (
      .rvfi_if    (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
      .support_if (support_logic_module_o_if.slave_mp),
      .*
    );


  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_data_independent_timing_assert #(
        .SECURE  (SECURE)
      ) xsecure_data_independent_timing_assert_i   (

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        //Interfaces:
        .rvfi_if    (rvfi_instr_if),
        .rvfi_cpuctrl (rvfi_csr_cpuctrl_if),

        //CSRs:
        .dataindtiming_enabled (core_i.xsecure_ctrl.cpuctrl.dataindtiming)
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_hardened_pc_assert #(
        .SECURE  (SECURE)
      ) xsecure_hardened_pc_assert_i   (

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        //CSRs:
        .pc_hardening_enabled (core_i.xsecure_ctrl.cpuctrl.pc_hardening),
        .dataindtiming_enabled (core_i.xsecure_ctrl.cpuctrl.dataindtiming),

        //Alert:
        .alert_major_due_to_pc_err (core_i.alert_i.pc_err_i),

        //IF:
        .if_valid (core_i.if_valid),
        .ptr_in_if (core_i.if_stage_i.ptr_in_if_o),
        .if_instr_cmpr (core_i.if_stage_i.compressed_decoder_i.is_compressed_o),
        .if_pc (core_i.pc_if),
        .dummy_insert (dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.dummy_insert),

        //ID:
        .id_ready (core_i.id_ready),
        .id_pc (core_i.id_stage_i.if_id_pipe_i.pc),
        .id_last_op (core_i.if_id_pipe.last_op),
        .id_first_op (core_i.if_id_pipe.first_op),
        .jump_in_id (core_i.controller_i.controller_fsm_i.jump_in_id),
        .kill_id (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.kill_id),
        .halt_id (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.halt_id),

        //EX:
        .ex_first_op (core_i.id_ex_pipe.first_op),
        .branch_in_ex (core_i.controller_i.controller_fsm_i.branch_in_ex),
        .kill_ex (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.kill_ex),
        .halt_ex (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.halt_ex),

        //Controll signals:
        .pc_set (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.pc_set),
        .pc_mux (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.pc_mux),

        //Signals to glitch check:
        .branch_target (core_i.ex_stage_i.branch_target_o),
        .branch_decision (core_i.ex_stage_i.alu_i.cmp_result_o),
        .jump_target (core_i.jump_target_id),
        .mepc (core_i.cs_registers_i.mepc_rdata)

      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_reduced_profiling_infrastructure_assert #(
        .SECURE  (SECURE)
      ) xsecure_reduced_profiling_infrastructure_assert_i   (

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        .mhpmevent (core_i.cs_registers_i.mhpmevent_rdata),
        .mhpmcounter (core_i.cs_registers_i.mhpmcounter_rdata),
        .mcountinhibit (core_i.cs_registers_i.mcountinhibit_rdata)
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_hardened_csrs_assert #(
        .SECURE  (SECURE)
      ) xsecure_hardened_csrs_assert_i   (

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        //Alert:
        .alert_major (core_i.alert_major_o),

        //CSRs:
        .mstateen0            (core_i.cs_registers_i.mstateen0_csr_i.rdata_q),
        .priv_lvl             (core_i.cs_registers_i.privlvl_user.priv_lvl_i.rdata_q),
        .jvt                  (core_i.cs_registers_i.jvt_csr_i.rdata_q),
        .mstatus              (core_i.cs_registers_i.mstatus_csr_i.rdata_q),
        .cpuctrl              (core_i.cs_registers_i.xsecure.cpuctrl_csr_i.rdata_q),
        .dcsr                 (core_i.cs_registers_i.gen_debug_csr.dcsr_csr_i.rdata_q),
        .mepc                 (core_i.cs_registers_i.mepc_csr_i.rdata_q),
        .mscratch             (core_i.cs_registers_i.mscratch_csr_i.rdata_q),

        //Shadows:
        .mstateen0_shadow     (core_i.cs_registers_i.mstateen0_csr_i.gen_hardened.shadow_q),
        .priv_lvl_shadow      (core_i.cs_registers_i.privlvl_user.priv_lvl_i.gen_hardened.shadow_q),
        .jvt_shadow           (core_i.cs_registers_i.jvt_csr_i.gen_hardened.shadow_q),
        .mstatus_shadow       (core_i.cs_registers_i.mstatus_csr_i.gen_hardened.shadow_q),
        .cpuctrl_shadow       (core_i.cs_registers_i.xsecure.cpuctrl_csr_i.gen_hardened.shadow_q),
        .dcsr_shadow          (core_i.cs_registers_i.gen_debug_csr.dcsr_csr_i.gen_hardened.shadow_q),
        .mepc_shadow          (core_i.cs_registers_i.mepc_csr_i.gen_hardened.shadow_q),
        .mscratch_shadow      (core_i.cs_registers_i.mscratch_csr_i.gen_hardened.shadow_q)

      );
  `endif

  if (CORE_PARAM_CLIC == 1) begin: gen_hardened_csrs_clic_assert
    `ifndef  COREV_ASSERT_OFF
      bind cv32e40s_wrapper
        uvmt_cv32e40s_xsecure_hardened_csrs_clic_assert #(
          .SECURE  (SECURE)
        ) xsecure_hardened_csrs_clic_assert_i   (

          //Signals:
          .clk_i      (clknrst_if.clk),
          .rst_ni     (clknrst_if.reset_n),

          //Alert:
          .alert_major (core_i.alert_major_o),

          //CSRs:
          .mcause             (core_i.cs_registers_i.clic_csrs.mcause_csr_i.rdata_q),
          .mtvt               (core_i.cs_registers_i.clic_csrs.mtvt_csr_i.rdata_q),
          .mtvec              (core_i.cs_registers_i.clic_csrs.mtvec_csr_i.rdata_q),
          .mintstatus         (core_i.cs_registers_i.clic_csrs.mintstatus_csr_i.rdata_q),
          .mintthresh         (core_i.cs_registers_i.clic_csrs.mintthresh_csr_i.rdata_q),

          //Shadows:
          .mcause_shadow      (core_i.cs_registers_i.clic_csrs.mcause_csr_i.gen_hardened.shadow_q),
          .mtvt_shadow        (core_i.cs_registers_i.clic_csrs.mtvt_csr_i.gen_hardened.shadow_q),
          .mtvec_shadow       (core_i.cs_registers_i.clic_csrs.mtvec_csr_i.gen_hardened.shadow_q),
          .mintstatus_shadow  (core_i.cs_registers_i.clic_csrs.mintstatus_csr_i.gen_hardened.shadow_q),
          .mintthresh_shadow  (core_i.cs_registers_i.clic_csrs.mintthresh_csr_i.gen_hardened.shadow_q)

        );
    `endif
  end : gen_hardened_csrs_clic_assert

  if (CORE_PARAM_CLIC == 0) begin: gen_hardened_csrs_interrupt_assert
    `ifndef  COREV_ASSERT_OFF
      bind cv32e40s_wrapper
        uvmt_cv32e40s_xsecure_hardened_csrs_interrupt_assert #(
          .SECURE  (SECURE)
        ) xsecure_hardened_csrs_interrupt_assert_i   (

          //Signals:
          .clk_i      (clknrst_if.clk),
          .rst_ni     (clknrst_if.reset_n),

          //Alert:
          .alert_major (core_i.alert_major_o),

          //CSRs:
          .mcause             (core_i.cs_registers_i.basic_mode_csrs.mcause_csr_i.rdata_q),
          .mtvec              (core_i.cs_registers_i.basic_mode_csrs.mtvec_csr_i.rdata_q),
          .mie                (core_i.cs_registers_i.basic_mode_csrs.mie_csr_i.rdata_q),

          //Shadows:
          .mcause_shadow      (core_i.cs_registers_i.basic_mode_csrs.mcause_csr_i.gen_hardened.shadow_q),
          .mtvec_shadow       (core_i.cs_registers_i.basic_mode_csrs.mtvec_csr_i.gen_hardened.shadow_q),
          .mie_shadow         (core_i.cs_registers_i.basic_mode_csrs.mie_csr_i.gen_hardened.shadow_q)
        );
    `endif
  end : gen_hardened_csrs_interrupt_assert



  if (CORE_PARAM_PMP_NUM_REGIONS > 0) begin: gen_hardened_csrs_pmp_assert
    localparam PMP_ADDR_WIDTH = (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_GRANULARITY > 0) ? 33 - uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_GRANULARITY : 32;

    pmpncfg_t pmpncfg[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_NUM_REGIONS];
    logic [PMP_ADDR_WIDTH-1:0] pmp_addr[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_NUM_REGIONS];

    logic [$bits(pmpncfg_t)-1:0] pmpncfg_shadow[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_NUM_REGIONS];
    logic [PMP_ADDR_WIDTH-1:0] pmp_addr_shadow[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_NUM_REGIONS];

    for (genvar n = 0; n < uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_NUM_REGIONS; n++) begin
      assign pmpncfg[n] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.csr_pmp.gen_pmp_csr[n].pmp_region.pmpncfg_csr_i.rdata_q;
      assign pmp_addr[n] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.csr_pmp.gen_pmp_csr[n].pmp_region.pmp_addr_csr_i.rdata_q;

      assign pmpncfg_shadow[n] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.csr_pmp.gen_pmp_csr[n].pmp_region.pmpncfg_csr_i.gen_hardened.shadow_q;
      assign pmp_addr_shadow[n] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.csr_pmp.gen_pmp_csr[n].pmp_region.pmp_addr_csr_i.gen_hardened.shadow_q;
    end


    `ifndef  COREV_ASSERT_OFF
      bind cv32e40s_wrapper
        uvmt_cv32e40s_xsecure_hardened_csrs_pmp_assert #(
          .SECURE  (SECURE),
          .PMP_ADDR_WIDTH (core_i.cs_registers_i.PMP_ADDR_WIDTH),
          .PMP_NUM_REGIONS (PMP_NUM_REGIONS)
        ) xsecure_hardened_csrs_pmp_assert_i   (

          //Signals:
          .clk_i      (clknrst_if.clk),
          .rst_ni     (clknrst_if.reset_n),

          //Alert:
          .alert_major (core_i.alert_major_o),

          //CSRs:
          .pmp_mseccfg        (core_i.cs_registers_i.csr_pmp.pmp_mseccfg_csr_i.rdata_q),
          .pmpncfg            (uvmt_cv32e40s_tb.gen_hardened_csrs_pmp_assert.pmpncfg),
          .pmp_addr           (uvmt_cv32e40s_tb.gen_hardened_csrs_pmp_assert.pmp_addr),

          //Shadows:
          .pmp_mseccfg_shadow (core_i.cs_registers_i.csr_pmp.pmp_mseccfg_csr_i.gen_hardened.shadow_q),
          .pmpncfg_shadow     (uvmt_cv32e40s_tb.gen_hardened_csrs_pmp_assert.pmpncfg_shadow),
          .pmp_addr_shadow    (uvmt_cv32e40s_tb.gen_hardened_csrs_pmp_assert.pmp_addr_shadow)
        );
    `endif

  end : gen_hardened_csrs_pmp_assert

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_register_file_ecc_assert #(
	    .SECURE	(SECURE)
      ) xsecure_register_file_ecc_assert_i 	(

        //Interfaces:
        .rvfi_if	  (rvfi_instr_if),

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        //Alert:
        .alert_major (core_i.alert_major_o),

        //Register file memory:
        .gpr_mem (core_i.register_file_wrapper_i.register_file_i.mem_gated),

        //Soruce registers:
        .rs1 (core_i.if_id_pipe.instr.bus_resp.rdata[19:15]),
        .rs2 (core_i.if_id_pipe.instr.bus_resp.rdata[24:20]),

        //Writing of GPRs:
        .gpr_we (core_i.rf_we_wb),
        .gpr_waddr (core_i.rf_waddr_wb),
        .gpr_wdata (core_i.rf_wdata_wb)

      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_security_alerts_assert #(
	    .SECURE	(SECURE)
      ) xsecure_security_alerts_assert_i 	(

        //Interfaces:
        .rvfi_if	  (rvfi_instr_if),
        .support_if (support_logic_module_o_if.slave_mp),

        //Signals:
        .rst_ni     (clknrst_if.reset_n),
        .clk_i      (clknrst_if.clk),

        //alerts:
        .alert_minor (core_i.alert_minor_o),
        .alert_major (core_i.alert_major_o),

        //wb:
        .wb_valid (core_i.wb_valid),
        .exception_in_wb (core_i.controller_i.controller_fsm_i.exception_in_wb),
        .exception_cause_wb (core_i.controller_i.controller_fsm_i.exception_cause_wb),

        //dummy and hint:
        .dummy_en (core_i.xsecure_ctrl.cpuctrl.rnddummy),
        .hint_en (core_i.xsecure_ctrl.cpuctrl.rndhint),
        .lfsr0_clock_en (core_i.cs_registers_i.xsecure.lfsr0_i.clock_en),
        .lfsr1_clock_en (core_i.cs_registers_i.xsecure.lfsr1_i.clock_en),
        .lfsr2_clock_en (core_i.cs_registers_i.xsecure.lfsr2_i.clock_en),
        .seed0_we       (core_i.cs_registers_i.xsecure.lfsr0_i.seed_we_i),
        .seed1_we       (core_i.cs_registers_i.xsecure.lfsr1_i.seed_we_i),
        .seed2_we       (core_i.cs_registers_i.xsecure.lfsr2_i.seed_we_i),
        .seed0_i        (core_i.cs_registers_i.xsecure.lfsr0_i.seed_i),
        .seed1_i        (core_i.cs_registers_i.xsecure.lfsr1_i.seed_i),
        .seed2_i        (core_i.cs_registers_i.xsecure.lfsr2_i.seed_i),
        .lfsr0_n        (core_i.cs_registers_i.xsecure.lfsr0_i.lfsr_n),
        .lfsr1_n        (core_i.cs_registers_i.xsecure.lfsr1_i.lfsr_n),
        .lfsr2_n        (core_i.cs_registers_i.xsecure.lfsr2_i.lfsr_n),

        //OBI:
        .obi_data_rvalid (core_i.data_rvalid_i),
        .obi_data_err (core_i.data_err_i),

        //NMI:
        .nmip (core_i.dcsr.nmip),

        //debug:
        .debug_mode (core_i.controller_i.controller_fsm_i.debug_mode_q)

      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_bus_protocol_hardening_assert #(
	    .SECURE	(SECURE)
      ) xsecure_bus_protocol_hardening_assert_i 	(

        //Interfaces:
        .support_if (support_logic_module_o_if.slave_mp),

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        //Alerts:
        .alert_major (core_i.alert_major_o),
        .bus_protocol_hardening_glitch (core_i.alert_i.itf_prot_err_i),

        //OBI:
        .obi_data_rvalid (core_i.m_c_obi_data_if.s_rvalid.rvalid),
        .obi_instr_rvalid (core_i.m_c_obi_instr_if.s_rvalid.rvalid),

        //Resp valids:
        .instr_if_mpu_resp (core_i.if_stage_i.prefetch_resp_valid),
        .lsu_mpu_resp (core_i.load_store_unit_i.resp_valid),

        //Counters:
        .lsu_rf_core_side_cnt (core_i.load_store_unit_i.response_filter_i.core_cnt_q),
        .lsu_rf_bus_side_cnt (core_i.load_store_unit_i.response_filter_i.bus_cnt_q)

      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_interface_integrity_assert #(
	    .SECURE	(SECURE),
        .ALBUF_DEPTH (core_i.if_stage_i.ALBUF_DEPTH),
        .ALBUF_CNT_WIDTH (core_i.if_stage_i.ALBUF_CNT_WIDTH)
      ) xsecure_interface_integrity_assert_i 	(

        //Interfaces:
        .support_if (support_logic_module_o_if.slave_mp),

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        //Alert:
        .alert_major (core_i.alert_major_o),
        .alert_major_due_to_integrity_err (core_i.alert_i.itf_int_err_i),

        //CSRs:
        .integrity_enabled (core_i.xsecure_ctrl.cpuctrl.integrity),
        .nmip (core_i.cs_registers_i.dcsr_rdata.nmip),
        .mcause_exception_code (core_i.cs_registers_i.mcause_rdata.exception_code),

        //OBI data:
        .obi_data_req_packet (core_i.m_c_obi_data_if.req_payload),
        .obi_data_resp_packet (core_i.m_c_obi_data_if.resp_payload),
        .obi_data_addr (core_i.data_addr_o),
        .obi_data_req (core_i.m_c_obi_data_if.s_req.req),
        .obi_data_reqpar (core_i.m_c_obi_data_if.s_req.reqpar),
        .obi_data_gnt (core_i.m_c_obi_data_if.s_gnt.gnt),
        .obi_data_gntpar (core_i.m_c_obi_data_if.s_gnt.gntpar),
        .obi_data_rvalid (core_i.m_c_obi_data_if.s_rvalid.rvalid),
        .obi_data_rvalidpar (core_i.m_c_obi_data_if.s_rvalid.rvalidpar),

        //OBI instr:
        .obi_instr_req_packet (core_i.m_c_obi_instr_if.req_payload),
        .obi_instr_resp_packet (core_i.m_c_obi_instr_if.resp_payload),
        .obi_instr_addr (core_i.instr_addr_o),
        .obi_instr_req (core_i.m_c_obi_instr_if.s_req.req),
        .obi_instr_reqpar (core_i.m_c_obi_instr_if.s_req.reqpar),
        .obi_instr_gnt (core_i.m_c_obi_instr_if.s_gnt.gnt),
        .obi_instr_gntpar (core_i.m_c_obi_instr_if.s_gnt.gntpar),
        .obi_instr_rvalid (core_i.m_c_obi_instr_if.s_rvalid.rvalid),
        .obi_instr_rvalidpar (core_i.m_c_obi_instr_if.s_rvalid.rvalidpar),

        //Register file memory:
        .gpr_mem (core_i.register_file_wrapper_i.register_file_i.mem_gated),
        .rf_we (core_i.rf_we_wb),
        .rf_waddr (core_i.rf_waddr_wb),
        .rf_wdata (core_i.rf_wdata_wb),

        //Alignment buffer:
        .alb_resp_i (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.resp_i),
        .alb_resp_q (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.resp_q),
        .alb_valid (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.valid_q),
        .alb_wptr (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.wptr),
        .alb_rptr1 (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.rptr),
        .alb_rptr2 (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.rptr2),

        //If:
        .if_valid (core_i.if_valid),
        .if_instr_integrity_err (core_i.if_stage_i.bus_resp.integrity_err),
        .if_instr_cmpr (core_i.if_stage_i.compressed_decoder_i.is_compressed_o),
        .if_instr_pc (core_i.if_stage_i.pc_if_o),
        .dummy_insert (dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.dummy_insert),

        //Id:
        .id_ready (core_i.id_ready),
        .id_instr_integrity_err (core_i.if_id_pipe.instr.bus_resp.integrity_err),
        .id_abort_op (dut_wrap.cv32e40s_wrapper_i.core_i.if_id_pipe.abort_op),
        .id_illegal_insn (dut_wrap.cv32e40s_wrapper_i.core_i.if_id_pipe.illegal_c_insn),

        //Wb:
        .wb_valid (core_i.wb_valid),
        .wb_integrity_err (core_i.ex_wb_pipe.instr.bus_resp.integrity_err),
        .wb_instr_opcode (core_i.ex_wb_pipe.instr.bus_resp.rdata[6:0]),
        .wb_exception (core_i.controller_i.controller_fsm_i.exception_in_wb),
        .wb_exception_code (core_i.controller_i.controller_fsm_i.exception_cause_wb),
        .data_integrity_err (core_i.load_store_unit_i.bus_resp.integrity_err),

        //MISC:
        .ctrl_fsm_cs (core_i.controller_i.controller_fsm_i.ctrl_fsm_cs),
        .pc_mux (dut_wrap.cv32e40s_wrapper_i.core_i.ctrl_fsm.pc_mux),
        .pc_set (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.ctrl_fsm_i.pc_set),
        .seq_valid (core_i.if_stage_i.seq_valid),
        .kill_if (core_i.ctrl_fsm.kill_if),
        .n_flush_q (core_i.if_stage_i.prefetch_unit_i.alignment_buffer_i.n_flush_q),
        .rchk_err_instr (core_i.if_stage_i.instruction_obi_i.rchk_err_resp),
        .rchk_err_data (core_i.load_store_unit_i.data_obi_i.rchk_err_resp)

      );
  `endif


  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_xsecure_dummy_and_hint_assert #(
	    .SECURE	(SECURE)
      ) xsecure_dummy_and_hint_assert_i 	(

        //Interfaces:
        .rvfi_if	  (rvfi_instr_if),
        .rvfi_mcountinhibit_if (rvfi_csr_mcountinhibit_if),
        .rvfi_dcsr_if (rvfi_csr_dcsr_if),

        //Signals:
        .clk_i      (clknrst_if.clk),
        .rst_ni     (clknrst_if.reset_n),

        .gated_clk_enabled (core_i.sleep_unit_i.clock_en),

        //CSRs:
        .rnddummy_enabled (core_i.xsecure_ctrl.cpuctrl.rnddummy),
        .rndhint_enabled (core_i.xsecure_ctrl.cpuctrl.rndhint),
        .dummy_freq (core_i.xsecure_ctrl.cpuctrl.rnddummyfreq),
        .mhpmcounter (core_i.cs_registers_i.mhpmcounter_rdata),
        .mcountinhibit (core_i.cs_registers_i.mcountinhibit_rdata),
        .csr_waddr(core_i.cs_registers_i.csr_waddr),

        //LFSR:
        .lfsr0_seed_we (core_i.cs_registers_i.xsecure.lfsr0_i.seed_we_i),
        .lfsr1_seed_we (core_i.cs_registers_i.xsecure.lfsr1_i.seed_we_i),
        .lfsr2_seed_we (core_i.cs_registers_i.xsecure.lfsr2_i.seed_we_i),
        .lfsr0_seed (core_i.cs_registers_i.xsecure.lfsr0_i.seed_i),
        .lfsr1_seed (core_i.cs_registers_i.xsecure.lfsr1_i.seed_i),
        .lfsr2_seed (core_i.cs_registers_i.xsecure.lfsr2_i.seed_i),
        .lfsr0 (core_i.cs_registers_i.xsecure.lfsr0_i.lfsr_q),
        .lfsr1 (core_i.cs_registers_i.xsecure.lfsr1_i.lfsr_q),
        .lfsr2 (core_i.cs_registers_i.xsecure.lfsr2_i.lfsr_q),
        .lfsr0_n (core_i.cs_registers_i.xsecure.lfsr0_i.lfsr_n),
        .lfsr1_n (core_i.cs_registers_i.xsecure.lfsr1_i.lfsr_n),
        .lfsr2_n (core_i.cs_registers_i.xsecure.lfsr2_i.lfsr_n),
        .lfsr0_clk_en (core_i.cs_registers_i.xsecure.lfsr0_i.clock_en),
        .lfsr1_clk_en (core_i.cs_registers_i.xsecure.lfsr1_i.clock_en),
        .lfsr2_clk_en (core_i.cs_registers_i.xsecure.lfsr2_i.clock_en),

        //IF:
        .if_hint  (core_i.if_stage_i.instr_hint),
        .if_dummy (core_i.if_stage_i.dummy_insert),
        .kill_if  (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.kill_if),
        .if_valid (core_i.if_valid),
        .ptr_in_if (core_i.if_stage_i.ptr_in_if_o),
        .if_first_op (core_i.if_stage_i.first_op),

        //ID:
        .operand_a (core_i.id_stage_i.operand_a),
        .operand_b (core_i.id_stage_i.operand_b),
        .id_instr (core_i.if_id_pipe.instr.bus_resp.rdata),
        .id_dummy (core_i.if_id_pipe.instr_meta.dummy),
        .id_hint (core_i.if_id_pipe.instr_meta.hint),
        .kill_id (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.kill_id),
        .id_ready (core_i.id_ready),
        .id_valid (core_i.id_valid),
        .id_last_op (core_i.id_stage_i.last_op),

        //EX:
        .kill_ex (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.kill_ex),
        .ex_ready (core_i.ex_ready),

        //WB:
        .kill_wb (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.kill_wb),
        .wb_dummy (core_i.ex_wb_pipe.instr_meta.dummy),
        .wb_hint (core_i.ex_wb_pipe.instr_meta.hint),
        .wb_valid (core_i.wb_valid),
        .wb_instr (core_i.ex_wb_pipe.instr.bus_resp.rdata),

        //Controller:
        .debug_mode (core_i.controller_i.controller_fsm_i.debug_mode_q),
        .stopcount_in_debug (core_i.cs_registers_i.debug_stopcount)
      );
  `endif


  // Debug assertion and coverage interface

  // Instantiate debug assertions

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper
      uvmt_cv32e40s_debug_cov_assert_if_t  debug_cov_assert_if (
        .id_valid               (core_i.id_stage_i.id_valid_o),
        .sys_fence_insn_i       (core_i.id_stage_i.decoder_i.sys_fencei_insn_o),

        .ex_stage_csr_en        (core_i.id_ex_pipe.csr_en),
        .ex_valid               (core_i.ex_stage_i.instr_valid),
        .ex_stage_instr_rdata_i (core_i.id_ex_pipe.instr.bus_resp.rdata),
        .ex_stage_pc            (core_i.id_ex_pipe.pc),

        .wb_stage_instr_rdata_i (core_i.ex_wb_pipe.instr.bus_resp.rdata),
        .wb_stage_instr_valid_i (core_i.ex_wb_pipe.instr_valid),
        .wb_stage_pc            (core_i.wb_stage_i.ex_wb_pipe_i.pc),
        .wb_err                 (core_i.ex_wb_pipe.instr.bus_resp.err),
        .wb_illegal             (core_i.ex_wb_pipe.illegal_insn),
        .wb_valid               (core_i.wb_stage_i.wb_valid_o),
        .wb_mpu_status          (core_i.ex_wb_pipe.instr.mpu_status),
        .illegal_insn_i         (core_i.ex_wb_pipe.illegal_insn),
        .sys_en_i               (core_i.ex_wb_pipe.sys_en),
        .sys_ecall_insn_i       (core_i.ex_wb_pipe.sys_ecall_insn),

        .ctrl_fsm_cs            (core_i.controller_i.controller_fsm_i.ctrl_fsm_cs),
        .debug_req_i            (core_i.controller_i.controller_fsm_i.debug_req_i),
        .debug_havereset        (core_i.debug_havereset_o),
        .debug_running          (core_i.debug_running_o),
        .debug_halted           (core_i.debug_halted_o),
        .debug_pc_o             (core_i.debug_pc_o),
        .debug_pc_valid_o       (core_i.debug_pc_valid_o),

        .ctrl_fsm_async_debug_allowed  (core_i.controller_i.controller_fsm_i.async_debug_allowed),
        .pending_sync_debug     (core_i.controller_i.controller_fsm_i.pending_sync_debug),
        .pending_async_debug    (core_i.controller_i.controller_fsm_i.pending_async_debug),
        .pending_nmi            (core_i.controller_i.controller_fsm_i.pending_nmi),
        .nmi_allowed            (core_i.controller_i.controller_fsm_i.nmi_allowed),
        .debug_mode_q           (core_i.controller_i.controller_fsm_i.debug_mode_q),
        .debug_mode_if          (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.debug_mode_if),
        .ctrl_halt_ex           (core_i.controller_i.controller_fsm_i.ctrl_fsm_o.halt_ex),
        .trigger_match_in_wb    (core_i.controller_i.controller_fsm_i.trigger_match_in_wb),
        .etrigger_in_wb         (core_i.controller_i.controller_fsm_i.etrigger_in_wb),
        .branch_in_ex           (core_i.controller_i.controller_fsm_i.branch_in_ex),

        .mie_q                  (core_i.cs_registers_i.mie_q),
        .dcsr_q                 (core_i.cs_registers_i.dcsr_q),
        .dpc_q                  (core_i.cs_registers_i.dpc_q),
        .dpc_n                  (core_i.cs_registers_i.dpc_n),
        .mcause_q               (core_i.cs_registers_i.mcause_q),
        .mtvec                  (core_i.cs_registers_i.mtvec_q),
        .mepc_q                 (core_i.cs_registers_i.mepc_q),
        .tdata1                 (core_i.cs_registers_i.tdata1_rdata),
        .tdata2                 (core_i.cs_registers_i.tdata2_rdata),
        .mcountinhibit_q        (core_i.cs_registers_i.mcountinhibit_q),
        .mcycle                 (core_i.cs_registers_i.mhpmcounter_q[0]),
        .minstret               (core_i.cs_registers_i.mhpmcounter_q[2]),
        .csr_we_int             (core_i.cs_registers_i.csr_we_int),

        // TODO: review this change from CV32E40S_HASH f6196bf to a26b194. It should be logically equivalent.
        //assign debug_cov_assert_if.inst_ret = core_i.cs_registers_i.inst_ret;
      // First attempt: this causes unexpected failures of a_minstret_count
      //assign debug_cov_assert_if.inst_ret = (core_i.id_valid &
      //                                       core_i.is_decoding);
      // Second attempt: (based on OK input).  This passes, but maybe only because p_minstret_count
      //                                       is the only property sensitive to inst_ret. Will
      //                                       this work in the general case?
      .inst_ret               (core_i.ctrl_fsm.mhpmevent.minstret),
      .csr_access             (core_i.ex_wb_pipe.csr_en),
      .csr_op                 (core_i.ex_wb_pipe.csr_op),
      .csr_addr               (core_i.ex_wb_pipe.csr_addr),
      .irq_ack_o              (core_i.irq_ack),
      .irq_id_o               (core_i.irq_id),
      .dm_halt_addr_i         (core_i.dm_halt_addr_i),
      .dm_exception_addr_i    (core_i.dm_exception_addr_i),
      .core_sleep_o           (core_i.core_sleep_o),
      .irq_i                  (core_i.irq_i),
      .pc_set                 (core_i.ctrl_fsm.pc_set),
      .boot_addr_i            (core_i.boot_addr_i),

      .is_wfi                 (),
      .dpc_will_hit           (),
      .addr_match             (),
      .is_ebreak              (),
      .is_cebreak             (),
      .is_dret                (),
      .is_mulhsu              (),
      .pending_enabled_irq    (),

      .*
    );
  `endif


    logic [31:0] tdata1_array[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DBG_NUM_TRIGGERS+1];
    logic [31:0] tdata2_array[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DBG_NUM_TRIGGERS+1];

    if (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DBG_NUM_TRIGGERS > 0) begin
      for (genvar t = 0; t < uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DBG_NUM_TRIGGERS; t++) begin
        assign tdata1_array[t] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.debug_triggers_i.gen_triggers.tdata1_rdata[t];
        assign tdata2_array[t] = dut_wrap.cv32e40s_wrapper_i.core_i.cs_registers_i.debug_triggers_i.gen_triggers.tdata2_rdata[t];
      end
      assign tdata1_array[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DBG_NUM_TRIGGERS] = '0;
      assign tdata2_array[uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DBG_NUM_TRIGGERS] = '0;

    end else begin
      assign tdata1_array = {'0};
      assign tdata2_array = {'0};
    end


  bind cv32e40s_wrapper
    uvmt_cv32e40s_support_logic_module_i_if_t support_logic_module_i_if (
      .clk     (core_i.clk),
      .rst_n (rst_ni),

      .if_instr (core_i.if_stage_i.prefetch_instr.bus_resp.rdata),
      .id_instr (core_i.if_id_pipe.instr.bus_resp.rdata),
      .ex_instr (core_i.id_ex_pipe.instr.bus_resp.rdata),
      .wb_instr (core_i.ex_wb_pipe.instr.bus_resp.rdata),

      .tdata1_array (uvmt_cv32e40s_tb.tdata1_array),
      .tdata2_array (uvmt_cv32e40s_tb.tdata2_array),

      .ctrl_fsm_o (core_i.controller_i.controller_fsm_i.ctrl_fsm_o),

      .fetch_enable        (core_i.fetch_enable),
      .debug_req_i         (core_i.debug_req_i),
      .irq_ack             (core_i.irq_ack),

      .wb_valid (core_i.wb_stage_i.wb_valid_o),
      .wb_tselect (core_i.cs_registers_i.tselect_rdata),
      .wb_tdata1 (core_i.cs_registers_i.tdata1_rdata),
      .wb_tdata2 (core_i.cs_registers_i.tdata2_rdata),

      .data_bus_rvalid (core_i.m_c_obi_data_if.s_rvalid.rvalid),
      .data_bus_req (core_i.m_c_obi_data_if.s_req.req),
      .data_bus_gnt (core_i.m_c_obi_data_if.s_gnt.gnt),
      .data_bus_gntpar (core_i.m_c_obi_data_if.s_gnt.gntpar),

      .instr_bus_rvalid (core_i.m_c_obi_instr_if.s_rvalid.rvalid),
      .instr_bus_req (core_i.m_c_obi_instr_if.s_req.req),
      .instr_bus_gnt (core_i.m_c_obi_instr_if.s_gnt.gnt),
      .instr_bus_gntpar (core_i.m_c_obi_instr_if.s_gnt.gntpar),

      //obi protocol between alignmentbuffer (ab) and instructoin (i) interface (i) mpu (m) is refered to as abiim
      .abiim_bus_rvalid (core_i.if_stage_i.prefetch_resp_valid),
      .abiim_bus_req (core_i.if_stage_i.prefetch_trans_ready),
      .abiim_bus_gnt (core_i.if_stage_i.prefetch_trans_valid),

      //obi protocol between LSU (l) mpu (m) and LSU (l) is refered to as lml
      .lml_bus_rvalid (core_i.load_store_unit_i.resp_valid),
      .lml_bus_req (core_i.load_store_unit_i.trans_ready),
      .lml_bus_gnt (core_i.load_store_unit_i.trans_valid),

      //obi protocol between LSU (l) respons (r) filter (f) and OBI (o) data (d) interface (i) is refered to as lrfodi
      .lrfodi_bus_rvalid (core_i.load_store_unit_i.bus_resp_valid),
      .lrfodi_bus_req (core_i.load_store_unit_i.buffer_trans_valid),
      .lrfodi_bus_gnt (core_i.load_store_unit_i.buffer_trans_ready),

      .req_instr_integrity (core_i.m_c_obi_instr_if.req_payload.integrity),
      .req_data_integrity (core_i.m_c_obi_data_if.req_payload.integrity)
  );

  bind cv32e40s_wrapper
    uvmt_cv32e40s_support_logic_module_o_if_t support_logic_module_o_if();

  `ifndef  COREV_ASSERT_OFF
    bind uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i.pmp.pmp_i
      uvmt_cv32e40s_pmp_assert#(
        .PMP_GRANULARITY  (PMP_GRANULARITY),
        .PMP_NUM_REGIONS  (PMP_NUM_REGIONS),
        .IS_INSTR_SIDE    (1'b1),
        .PMP_MSECCFG_RV   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_MSECCFG_RV)
      )
      u_pmp_assert_if_stage(.rst_n          (clknrst_if.reset_n),
                            .bus_trans_dbg  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i.bus_trans_o.dbg),
                            .obi_addr       (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_addr_o),
                            .obi_gnt        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_gnt_i),
                            .obi_req        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_req_o),
                            .rvfi_pc_rdata  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_pc_rdata),
                            .rvfi_valid     (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_valid),
                            .*);
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i.pmp.pmp_i
      uvmt_cv32e40s_pmp_assert#(
        .PMP_GRANULARITY  (PMP_GRANULARITY),
        .PMP_NUM_REGIONS  (PMP_NUM_REGIONS),
        .IS_INSTR_SIDE    (1'b0),
        .PMP_MSECCFG_RV   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_MSECCFG_RV)
      )
      u_pmp_assert_lsu(.rst_n          (clknrst_if.reset_n),
                       .bus_trans_dbg  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i.bus_trans_o.dbg),
                       .obi_addr       (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_addr_o),
                       .obi_gnt        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_gnt_i),
                       .obi_req        (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_req_o),
                       .rvfi_pc_rdata  (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_pc_rdata),
                       .rvfi_valid     (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_valid),
                       .*);
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.rvfi_i
      uvmt_cv32e40s_pmprvfi_assert #(
        .PMP_GRANULARITY (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_GRANULARITY),
        .PMP_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_NUM_REGIONS)
      ) pmprvfi_assert_i (
        .rvfi_if        (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
        .support_if     (support_logic_module_o_if.slave_mp),
        .rvfi_mem_addr  (rvfi_mem_addr [31:0]),
        .rvfi_mem_wmask (rvfi_mem_wmask[ 3:0]),
        .rvfi_mem_rmask (rvfi_mem_rmask[ 3:0]),
        .*
      );
  `endif


  // PMA Asserts & Covers

  wire pma_status_t  pma_status_instr;
  wire pma_status_t  pma_status_data;
  wire pma_status_t  pma_status_rvfidata_word0lowbyte;
  wire pma_status_t  pma_status_rvfidata_word0highbyte;

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i
      uvmt_cv32e40s_pma_model #(
        .DM_REGION_END   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (1'b 1),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG)
      ) pma_model_instr_i (
        .addr_i       (pma_i.trans_addr_i),
        .dbg          (core_trans_i.dbg),
        .jvt_q        (core_i.cs_registers_i.jvt_q),
        .pma_status_o (uvmt_cv32e40s_tb.pma_status_instr),
        .*
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i
      uvmt_cv32e40s_pma_model #(
        .DM_REGION_END   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (1'b 0),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG)
      ) pma_model_data_i (
        .addr_i       (pma_i.trans_addr_i),
        .dbg          (core_trans_i.dbg),
        .jvt_q        (core_i.cs_registers_i.jvt_q),
        .pma_status_o (uvmt_cv32e40s_tb.pma_status_data),
        .*
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i
      uvmt_cv32e40s_pma_model #(
        .DM_REGION_END   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (1'b 0),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG)
      ) pma_model_rvfidata_low_i (
        .clk                  (clknrst_if.clk),
        .rst_n                (clknrst_if.reset_n),
        .addr_i               (rvfi_instr_if.rvfi_mem_addr[31:0]),
        .core_trans_pushpop_i (rvfi_instr_if.is_pushpop),
        .dbg                  (rvfi_instr_if.rvfi_dbg_mode),
        .jvt_q                (rvfi_csr_jvt_if.rvfi_csr_rdata),
        .load_access          (|rvfi_instr_if.rvfi_mem_rmask),
        .misaligned_access_i  (rvfi_instr_if.is_split_datatrans_intended),
        .pma_status_o         (uvmt_cv32e40s_tb.pma_status_rvfidata_word0lowbyte)
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i
      uvmt_cv32e40s_pma_model #(
        .DM_REGION_END   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (1'b 0),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG)
      ) pma_model_rvfidata_high_i (
        .clk                  (clknrst_if.clk),
        .rst_n                (clknrst_if.reset_n),
        .addr_i               (rvfi_instr_if.rvfi_mem_addr_word0highbyte),
          // TODO:WARNING:silabs-robin Should use "instr_mem_addr_word0highbyte"?
        .core_trans_pushpop_i (rvfi_instr_if.is_pushpop),
        .dbg                  (rvfi_instr_if.rvfi_dbg_mode),
        .jvt_q                (rvfi_csr_jvt_if.rvfi_csr_rdata),
        .load_access          (|rvfi_instr_if.rvfi_mem_rmask),
        .misaligned_access_i  (rvfi_instr_if.is_split_datatrans_intended),
        .pma_status_o         (uvmt_cv32e40s_tb.pma_status_rvfidata_word0highbyte)
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i
      uvmt_cv32e40s_pma_assert #(
        .CORE_REQ_TYPE   (cv32e40s_pkg::obi_inst_req_t),
        .DM_REGION_END   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (1),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG)
      ) pma_assert_instr_i (
        .obi_memory_if    (dut_wrap.obi_instr_if),
        .rvfi_instr_if    (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
        .writebuf_ready_o ('0),
        .writebuf_trans_i ('0),
        .writebuf_trans_o ('0),
        .pma_status_i     (uvmt_cv32e40s_tb.pma_status_instr),
        .*
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i
      uvmt_cv32e40s_pma_assert #(
        .CORE_REQ_TYPE   (cv32e40s_pkg::obi_data_req_t),
        .DM_REGION_END   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_END),
        .DM_REGION_START (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_START),
        .IS_INSTR_SIDE   (0),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
        .PMA_CFG         (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG)
      ) pma_assert_data_i (
        .obi_memory_if    (dut_wrap.obi_data_if),
        .rvfi_instr_if    (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
        .writebuf_ready_o (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.ready_o),
        .writebuf_trans_i (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.trans_i),
        .writebuf_trans_o (dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.write_buffer_i.trans_o),
        .pma_status_i     (uvmt_cv32e40s_tb.pma_status_data),
        .*
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i
      uvmt_cv32e40s_pma_cov #(
        .CORE_REQ_TYPE   (cv32e40s_pkg::obi_inst_req_t),
        .IS_INSTR_SIDE   (1'b 1),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS)
      ) pma_cov_instr_i (
        .clk_ungated                         (clknrst_if.clk),
        .pma_status_i                        (uvmt_cv32e40s_tb.pma_status_instr),
        .pma_status_rvfidata_word0lowbyte_i  (uvmt_cv32e40s_tb.pma_status_rvfidata_word0lowbyte),
        .pma_status_rvfidata_word0highbyte_i (uvmt_cv32e40s_tb.pma_status_rvfidata_word0highbyte),
        .rvfi_if                             (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
        .*
      );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind  dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i
      uvmt_cv32e40s_pma_cov #(
        .CORE_REQ_TYPE   (cv32e40s_pkg::obi_data_req_t),
        .IS_INSTR_SIDE   (1'b 0),
        .PMA_NUM_REGIONS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS)
      ) pma_cov_data_i (
        .clk_ungated                         (clknrst_if.clk),
        .pma_status_i                        (uvmt_cv32e40s_tb.pma_status_data),
        .pma_status_rvfidata_word0lowbyte_i  (uvmt_cv32e40s_tb.pma_status_rvfidata_word0lowbyte),
        .pma_status_rvfidata_word0highbyte_i (uvmt_cv32e40s_tb.pma_status_rvfidata_word0highbyte),
        .rvfi_if                             (dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if),
        .*
      );
  `endif


  // Support Logic

  bind cv32e40s_wrapper uvmt_cv32e40s_support_logic u_support_logic(.rvfi (rvfi_instr_if),
                                                                    .in_support_if (support_logic_module_i_if.driver_mp),
                                                                    .out_support_if (support_logic_module_o_if.master_mp),
                                                                    .data_obi_if (dut_wrap.obi_data_if),
                                                                    .instr_obi_if (dut_wrap.obi_instr_if)
                                                                    );


  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper uvmt_cv32e40s_debug_assert u_debug_assert(.rvfi(rvfi_instr_if),
                                                                    .csr_dcsr(rvfi_csr_dcsr_if),
                                                                    .csr_dpc(rvfi_csr_dpc_if),
                                                                    .csr_dscratch0(rvfi_csr_dscratch0_if),
                                                                    .csr_dscratch1(rvfi_csr_dscratch1_if),
                                                                    .csr_mepc(rvfi_csr_mepc_if),
                                                                    .csr_mstatus(rvfi_csr_mstatus_if),
                                                                    .csr_mcause(rvfi_csr_mcause_if),
                                                                    .csr_mtvec(rvfi_csr_mtvec_if),
                                                                    .csr_tdata1(rvfi_csr_tdata1_if),
                                                                    .csr_tdata2(rvfi_csr_tdata2_if),
                                                                    .instr_obi(dut_wrap.obi_instr_if),
                                                                    .data_obi(dut_wrap.obi_data_if),
                                                                    .cov_assert_if(debug_cov_assert_if),
                                                                    .support_if (support_logic_module_o_if.slave_mp)
                                                                    );
  `endif

  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper uvmt_cv32e40s_triggers_assert_cov debug_trigger_assert_i(
      .tdata1_array (uvmt_cv32e40s_tb.tdata1_array),
      .priv_lvl (core_i.priv_lvl),
      .rvfi_if (rvfi_instr_if),
      .clknrst_if (dut_wrap.clknrst_if),
      .support_if (support_logic_module_o_if.slave_mp),
      .tdata1_if (rvfi_csr_tdata1_if),
      .tdata2_if (rvfi_csr_tdata2_if),
      .tinfo_if (rvfi_csr_tinfo_if),
      .tselect_if (rvfi_csr_tselect_if),
      .dcsr_if (rvfi_csr_dcsr_if),
      .dpc_if (rvfi_csr_dpc_if)
    );
  `endif


  `ifndef  COREV_ASSERT_OFF
    bind cv32e40s_wrapper uvmt_cv32e40s_zc_assert u_zc_assert(.rvfi(rvfi_instr_if),
                                                              .support_if(support_logic_module_o_if.slave_mp)
                                                              );
  `endif

  `ifndef  COREV_ASSERT_OFF
    `ifdef  PARAM_SET_0
      `include  "cvverif_sva_binds.svh"
    `endif
  `endif

    //uvmt_cv32e40s_rvvi_handcar u_rvvi_handcar();

    // IMPERAS DV
    `ifndef FORMAL
      //uvmt_cv32e40s_imperas_dv_wrap imperas_dv (rvvi_if);
      uvmt_cv32e40s_reference_model_wrap reference_model (rvvi_if);
    `endif

   /**
    * Test bench entry point.
    */
   `ifndef FORMAL // Formal ignores initial blocks, avoids unnecessary warning
   initial begin : test_bench_entry_point

     // Specify time format for simulation (units_number, precision_number, suffix_string, minimum_field_width)
     $timeformat(-9, 3, " ns", 8);

     //uvm_config_db#(virtual uvmt_imperas_dv_if_t)::set(.cntxt(null), .inst_name("uvm_test_top"), .field_name("idv_support_vif"), .value(imperas_dv_if));
     uvm_config_db#(virtual uvmt_reference_model_if_t)::set(.cntxt(null), .inst_name("uvm_test_top"), .field_name("rm_support_vif"), .value(reference_model_if));
     // Add interfaces handles to uvm_config_db
     uvm_config_db#(virtual uvma_debug_if_t             )::set(.cntxt(null), .inst_name("*.env.debug_agent"),            .field_name("vif"),           .value(debug_if));
     uvm_config_db#(virtual uvma_clknrst_if_t           )::set(.cntxt(null), .inst_name("*.env.clknrst_agent"),          .field_name("vif"),           .value(clknrst_if));
     uvm_config_db#(virtual uvma_interrupt_if_t         )::set(.cntxt(null), .inst_name("*.env.interrupt_agent"),        .field_name("vif"),           .value(interrupt_if));
     uvm_config_db#(virtual uvma_wfe_wu_if_t            )::set(.cntxt(null), .inst_name("*.env.wfe_wu_agent"),           .field_name("vif"),           .value(wfe_wu_if));
     uvm_config_db#(virtual uvma_clic_if_t#(
       .CLIC_ID_WIDTH(uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC_ID_WIDTH)
     ))::set(.cntxt(null), .inst_name("*.env.clic_agent"), .field_name("vif"), .value(clic_if));

     uvm_config_db#(virtual uvma_obi_memory_if_t#(
       .AUSER_WIDTH(ENV_PARAM_INSTR_AUSER_WIDTH),
       .WUSER_WIDTH(ENV_PARAM_INSTR_WUSER_WIDTH),
       .RUSER_WIDTH(ENV_PARAM_INSTR_RUSER_WIDTH),
       .ADDR_WIDTH(ENV_PARAM_INSTR_ADDR_WIDTH),
       .DATA_WIDTH(ENV_PARAM_INSTR_DATA_WIDTH),
       .ID_WIDTH(ENV_PARAM_INSTR_ID_WIDTH),
       .ACHK_WIDTH(ENV_PARAM_INSTR_ACHK_WIDTH),
       .RCHK_WIDTH(ENV_PARAM_INSTR_RCHK_WIDTH)
     ))::set(.cntxt(null), .inst_name("*.env.obi_memory_instr_agent"), .field_name("vif"), .value(obi_instr_if) );
     uvm_config_db#(virtual uvma_obi_memory_if_t#(
       .AUSER_WIDTH(ENV_PARAM_DATA_AUSER_WIDTH),
       .WUSER_WIDTH(ENV_PARAM_DATA_WUSER_WIDTH),
       .RUSER_WIDTH(ENV_PARAM_DATA_RUSER_WIDTH),
       .ADDR_WIDTH(ENV_PARAM_DATA_ADDR_WIDTH),
       .DATA_WIDTH(ENV_PARAM_DATA_DATA_WIDTH),
       .ID_WIDTH(ENV_PARAM_DATA_ID_WIDTH),
       .ACHK_WIDTH(ENV_PARAM_DATA_ACHK_WIDTH),
       .RCHK_WIDTH(ENV_PARAM_DATA_RCHK_WIDTH)
     ))::set(.cntxt(null), .inst_name("*.env.obi_memory_data_agent"),  .field_name("vif"), .value(obi_data_if) );
     uvm_config_db#(virtual uvma_fencei_if_t            )::set(.cntxt(null), .inst_name("*.env.fencei"),                 .field_name("vif"),           .value(fencei_if));
     uvm_config_db#(virtual uvma_rvfi_instr_if_t        )::set(.cntxt(null), .inst_name("*.env.rvfi_agent"),             .field_name("instr_vif0"),    .value(dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if));
     uvm_config_db#(virtual uvma_fencei_if_t            )::set(.cntxt(null), .inst_name("*.env.fencei_agent"),           .field_name("fencei_vif"),    .value(fencei_if)  );
     uvm_config_db#(virtual uvmt_cv32e40s_vp_status_if_t)::set(.cntxt(null), .inst_name("*"),                            .field_name("vp_status_vif"), .value(vp_status_if) );
     uvm_config_db#(virtual uvma_interrupt_if_t         )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("intr_vif"),      .value(interrupt_if) );
     uvm_config_db#(virtual uvma_debug_if_t             )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("debug_vif"),     .value(debug_if)     );
     uvm_config_db#(virtual uvma_wfe_wu_if_t            )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("wfe_wu_vif"),    .value(wfe_wu_if)     );
     uvm_config_db#(virtual uvma_clic_if_t#(
       .CLIC_ID_WIDTH(uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC_ID_WIDTH)
     ))::set(.cntxt(null), .inst_name("*.env"), .field_name("clic_vif"), .value(clic_if) );
//     uvm_config_db#(virtual uvmt_cv32e40s_debug_cov_assert_if_t)::set(.cntxt(null), .inst_name("*.env"),                 .field_name("debug_cov_vif"),    .value(debug_cov_assert_if));
     `RVFI_CSR_UVM_CONFIG_DB_SET(cpuctrl)
     `RVFI_CSR_UVM_CONFIG_DB_SET(jvt)
     `RVFI_CSR_UVM_CONFIG_DB_SET(marchid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcause)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcounteren)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcountinhibit)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcycle)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcycleh)
     `RVFI_CSR_UVM_CONFIG_DB_SET(menvcfg)
     `RVFI_CSR_UVM_CONFIG_DB_SET(menvcfgh)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mepc)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhartid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mie)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mimpid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(minstret)
     `RVFI_CSR_UVM_CONFIG_DB_SET(minstreth)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mip)
     `RVFI_CSR_UVM_CONFIG_DB_SET(misa)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mscratch)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen0h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen1h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen2h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstateen3h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstatus)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstatush)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mtval)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mtvec)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mvendorid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mseccfg)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mseccfgh)

     `RVFI_CSR_UVM_CONFIG_DB_SET(dcsr)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dpc)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dscratch0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dscratch1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tselect)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tinfo)

     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg15)

     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr31)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr32)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr33)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr34)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr35)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr36)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr37)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr38)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr39)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr40)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr41)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr42)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr43)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr44)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr45)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr46)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr47)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr48)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr49)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr50)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr51)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr52)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr53)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr54)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr55)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr56)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr57)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr58)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr59)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr60)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr61)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr62)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr63)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent31)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter31)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter3h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter4h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter5h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter6h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter7h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter8h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter9h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter10h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter11h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter12h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter13h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter14h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter15h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter16h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter17h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter18h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter19h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter20h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter21h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter22h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter23h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter24h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter25h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter26h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter27h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter28h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter29h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter30h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter31h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mconfigptr)

     `RVFI_CSR_UVM_CONFIG_DB_SET(secureseed0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(secureseed1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(secureseed2)

     `ifdef CLIC_EN
       // TODO:silabs-robin  What about when using "PARAM_SET_0"?
       `RVFI_CSR_UVM_CONFIG_DB_SET(mintstatus)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mintthresh)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mnxti)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mscratchcsw)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mscratchcswl)
       `RVFI_CSR_UVM_CONFIG_DB_SET(mtvt)
     `endif

     // IMPERAS_DV interface
     if ($test$plusargs("USE_ISS")) begin
       uvm_config_db#(virtual rvviTrace)::set(.cntxt(null), .inst_name("*.env.rvvi_agent"), .field_name("rvvi_vif"), .value(rvvi_if));
     end

     // Virtual Peripheral Status interface
     uvm_config_db#(virtual uvmt_cv32e40s_vp_status_if_t              )::set(.cntxt(null), .inst_name("*"), .field_name("vp_status_vif"),       .value(vp_status_if)      );
     uvm_config_db#(virtual uvme_cv32e40s_core_cntrl_if_t             )::set(.cntxt(null), .inst_name("*"), .field_name("core_cntrl_vif"),      .value(core_cntrl_if)     );
     uvm_config_db#(virtual uvmt_cv32e40s_debug_cov_assert_if_t       )::set(.cntxt(null), .inst_name("*.env"), .field_name("debug_cov_vif"),.value(dut_wrap.cv32e40s_wrapper_i.debug_cov_assert_if));
     uvm_config_db#(virtual uvmt_cv32e40s_support_logic_module_o_if_t )::set(.cntxt(null), .inst_name("*.env"), .field_name("support_logic_vif"),.value(dut_wrap.cv32e40s_wrapper_i.support_logic_module_o_if));

     // Make the DUT Wrapper Virtual Peripheral's status outputs available to the base_test
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("tp"),     .value(1'b0)        );
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("tf"),     .value(1'b0)        );
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("evalid"), .value(1'b0)        );
     uvm_config_db#(bit[31:0])::set(.cntxt(null), .inst_name("*"), .field_name("evalue"), .value(32'h00000000));

     // DUT and ENV parameters
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_INSTR_ADDR_WIDTH"),  .value(ENV_PARAM_INSTR_ADDR_WIDTH) );
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_INSTR_DATA_WIDTH"),  .value(ENV_PARAM_INSTR_DATA_WIDTH) );
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_RAM_ADDR_WIDTH"),    .value(ENV_PARAM_RAM_ADDR_WIDTH)   );

     // Run test
     uvm_top.enable_print_topology = 0; // ENV coders enable this as a debug aid
     uvm_top.finish_on_completion  = 1;
     uvm_top.run_test();
   end : test_bench_entry_point
   `endif

   assign core_cntrl_if.clk = clknrst_if.clk;

   // Capture the test status and exit pulse flags
   // TODO: put this logic in the vp_status_if (makes it easier to pass to ENV)
   `ifndef FORMAL  // uvm db not used in formal
     always @(posedge clknrst_if.clk) begin
       if (!clknrst_if.reset_n) begin
         tp     <= 1'b0;
         tf     <= 1'b0;
         evalid <= 1'b0;
         evalue <= 32'h00000000;
       end
       else begin
         if (vp_status_if.tests_passed) begin
           tp <= 1'b1;
           uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("tp"), .value(1'b1));
         end
         if (vp_status_if.tests_failed) begin
           tf <= 1'b1;
           uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("tf"), .value(1'b1));
         end
         if (vp_status_if.exit_valid) begin
           evalid <= 1'b1;
           uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("evalid"), .value(1'b1));
         end
         if (vp_status_if.exit_valid) begin
           evalue <= vp_status_if.exit_value;
           uvm_config_db#(bit[31:0])::set(.cntxt(null), .inst_name("*"), .field_name("evalue"), .value(vp_status_if.exit_value));
         end
       end
     end
   `endif  // FORMAL


   /**
    * End-of-test summary printout.
    */
   `ifndef FORMAL // Formal ignores final blocks, this avoids unnecessary warning
   final begin: end_of_test
      string             summary_string;
      uvm_report_server  rs;
      int                err_count;
      int                warning_count;
      int                fatal_count;
      static bit         sim_finished = 0;

      static string  red   = "\033[31m\033[1m";
      static string  green = "\033[32m\033[1m";
      static string  reset = "\033[0m";

      rs            = uvm_top.get_report_server();
      err_count     = rs.get_severity_count(UVM_ERROR);
      warning_count = rs.get_severity_count(UVM_WARNING);
      fatal_count   = rs.get_severity_count(UVM_FATAL);

      if ($test$plusargs("USE_ISS")) begin
         void'(rvviApiPkg::rvviRefShutdown());
      end

      void'(uvm_config_db#(bit)::get(null, "", "sim_finished", sim_finished));

      `uvm_info("DV_WRAP", $sformatf("\n%m: *** Test Summary ***\n"), UVM_DEBUG);

      if (sim_finished && (err_count == 0) && (fatal_count == 0)) begin
         $display("    PPPPPPP    AAAAAA    SSSSSS    SSSSSS   EEEEEEEE  DDDDDDD     ");
         $display("    PP    PP  AA    AA  SS    SS  SS    SS  EE        DD    DD    ");
         $display("    PP    PP  AA    AA  SS        SS        EE        DD    DD    ");
         $display("    PPPPPPP   AAAAAAAA   SSSSSS    SSSSSS   EEEEE     DD    DD    ");
         $display("    PP        AA    AA        SS        SS  EE        DD    DD    ");
         $display("    PP        AA    AA  SS    SS  SS    SS  EE        DD    DD    ");
         $display("    PP        AA    AA   SSSSSS    SSSSSS   EEEEEEEE  DDDDDDD     ");
         $display("    ----------------------------------------------------------");
         if (warning_count == 0) begin
           $display("                        SIMULATION PASSED                     ");
         end
         else begin
           $display("                 SIMULATION PASSED with WARNINGS              ");
         end
         $display("    ----------------------------------------------------------");
      end
      else begin
         $display("    FFFFFFFF   AAAAAA   IIIIII  LL        EEEEEEEE  DDDDDDD       ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FFFFF     AAAAAAAA    II    LL        EEEEE     DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA  IIIIII  LLLLLLLL  EEEEEEEE  DDDDDDD       ");

         if (sim_finished == 0) begin
            $display("    --------------------------------------------------------");
            $display("                   SIMULATION FAILED - ABORTED              ");
            $display("    --------------------------------------------------------");
         end
         else begin
            $display("    --------------------------------------------------------");
            $display("                       SIMULATION FAILED                    ");
            $display("    --------------------------------------------------------");
         end
      end
      // If there are any liveness assertions still pending at this time,
      // kill all of them to prevent false failures after end of test.
      // Actual failures _should_ have been caught and logged at this time
      // This is needed as the core is not necessarily terminated by software,
      // and there may be outstanding transactions.
      $assertkill();
   end
   `endif

endmodule : uvmt_cv32e40s_tb
`default_nettype wire

`endif // __UVMT_CV32E40S_TB_SV__
