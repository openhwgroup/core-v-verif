// ----------------------------------------------------------------------------
// Copyright 2023 CEA*
// *Commissariat a l'Energie Atomique et aux Energies Alternatives (CEA)
//
// SPDX-License-Identifier: Apache-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//    http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//[END OF HEADER]
// ----------------------------------------------------------------------------
// ----------------------------------------------------------------------------
// ----------------------------------------------------------------------------
// ----------------------------------------------------------------------------
//  Description : Package with defines for XRTL portion of clock IF
//                
// 
// ----------------------------------------------------------------------------

package clock_mon_vif_xrtl_pkg;

  class xrtl_clock_mon_vif_c;

    // ----------------------------------------------------------------------
    // Name
    // ----------------------------------------------------------------------

    protected string name;

    // ----------------------------------------------------------------------
    // Constructor
    // ----------------------------------------------------------------------

    function new( string name_in ) ;
        name = name_in;
    endfunction : new

  endclass : xrtl_clock_mon_vif_c

endpackage : clock_mon_vif_xrtl_pkg
