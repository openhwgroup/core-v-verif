// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


`ifndef __UVMA_DEBUG_IF_CHK_SV__
`define __UVMA_DEBUG_IF_CHK_SV__


/**
 * Encapsulates assertions targeting uvma_debug_if_t.
 */
module uvma_debug_if_chk(
   uvma_debug_if_t  debug_if
);

   `pragma protect begin

   // TODO Add assertions to uvma_debug_if_chk

   `pragma protect end

endmodule : uvma_debug_if_chk


`endif // __UVMA_DEBUG_IF_CHK_SV__
