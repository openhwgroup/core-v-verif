POST_INC_LOAD,
POST_INC_STORE,
EVENT_LOAD,
HWLOOP,
BITMANIP,
ALU,
BRANCH_IMM,
MAC,
SIMD,
