
// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// 
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     https://solderpad.org/licenses/
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 

// This file specifies all interfaces used by the CV32E40P test bench (uvmt_cv32e40p_tb).
// Most interfaces support tasks to allow control by the ENV or test cases.

`ifndef __UVMT_CV32E40P_TB_IFS_SV__
`define __UVMT_CV32E40P_TB_IFS_SV__


/**
 * clocks and reset
 */
interface uvmt_cv32e40p_clk_gen_if (output logic core_clock, output logic core_reset_n);

   import uvm_pkg::*;
   
   bit       start_clk               = 0;
   // TODO: get the uvme_cv32e40p_* values from random ENV CFG members.
   realtime  core_clock_period       = 1500ps; // uvme_cv32e40p_clk_period * 1ps;
   realtime  reset_deassert_duration = 7400ps; // uvme_cv32e40p_reset_deassert_duarion * 1ps;
   realtime  reset_assert_duration   = 7400ps; // uvme_cv32e40p_reset_assert_duarion * 1ps;
   
   
   /**
    * Generates clock and reset signals.
    * If reset_n comes up de-asserted (1'b1), wait a bit, then assert, then de-assert
    * Otherwise, leave reset asserted, wait a bit, then de-assert.
    */
   initial begin
      core_clock   = 0; // uvme_cv32e40p_clk_initial_value;
      core_reset_n = 0; // uvme_cv32e40p_reset_initial_value;
      wait (start_clk);
      fork
         forever begin
            #(core_clock_period/2) core_clock = ~core_clock;
         end
         begin
           if (core_reset_n == 1'b1) #(reset_deassert_duration);
           core_reset_n = 1'b0;
           #(reset_assert_duration);
           core_reset_n = 1'b1;
         end
      join_none
   end
   
   /**
    * Sets clock period in ps.
    */
   function static void set_clk_period ( real clk_period );
      core_clock_period = clk_period * 1ps;
   endfunction : set_clk_period
   
   /** Triggers the generation of clk. */
   function static void start();
      start_clk = 1;
      `uvm_info("CLK_GEN_IF", "uvmt_cv32e40p_clk_gen_if.start() called", UVM_NONE)
   endfunction : start
   
endinterface : uvmt_cv32e40p_clk_gen_if

/**
 * Status information generated by the Virtual Peripherals in the DUT WRAPPER memory.
 */
interface uvmt_cv32e40p_vp_status_if (
                                  output reg        tests_passed,
                                  output reg        tests_failed,
                                  output reg        exit_valid,
                                  output reg [31:0] exit_value
                                 );

  import uvm_pkg::*;

  // TODO: X/Z checks
  initial begin
  end

endinterface : uvmt_cv32e40p_vp_status_if



/**
 * Core status signals.
 */
interface uvmt_cv32e40p_core_status_if (
                                    input  wire        core_busy,
                                    input  logic       sec_lvl
                                   );

  import uvm_pkg::*;

endinterface : uvmt_cv32e40p_core_status_if

/**
 * ISA coverage interface
 * ISS wrapper will fill in ins (instruction) and fire ins_valid event
 */
interface uvmt_cv32e40p_isa_covg_if;

  import uvm_pkg::*;
  import uvme_cv32e40p_pkg::*;

  event ins_valid;
  ins_t ins;

endinterface : uvmt_cv32e40p_isa_covg_if

/**
 * Step and compare interface
 * Xcelium does not support event types in the module port list
 */
interface uvmt_cv32e40p_step_compare_if;

  import uvm_pkg::*;

  // From RTL riscv_tracer.sv
  typedef struct {
     logic [ 5:0] addr;
     logic [31:0] value;
   } reg_t;

   event        ovp_cpu_valid;      // Indicate instruction successfully retired
   event        ovp_cpu_trap;       // Indicate exception occured 
   event        ovp_cpu_halt;       // Indicate exception occured 
   bit   [31:0] ovp_cpu_PCr;        // Was iss_wrap.cpu.PCr
   logic [31:0] ovp_cpu_GPR[32];
   bit          ovp_cpu_state_idle;
   bit          ovp_cpu_state_stepi;
   bit          ovp_cpu_state_stop;
   bit          ovp_cpu_state_cont;

   event        riscv_retire;       // Was riscv_core.riscv_tracer_i.retire
   event        riscv_trap;         // new event to indicate RTL took a trap
   event        riscv_halt;         // new event to indicate RTL took a halt
   
   logic [31:0] insn_pc;
   logic [31:0][31:0] riscy_GPR;    // packed dimensions, register index by data width
   logic        deferint_prime;     // Stages deferint for the ISS deferint signal
   logic        deferint_prime_ack; // Set low if deferint_prime was set due to interrupt ack (as opposed to wakeup)

   int  num_pc_checks;
   int  num_gpr_checks;
   int  num_csr_checks;

   // Report on the checkers at the end of simulation
   function void report_step_compare();
      if (num_pc_checks > 0) begin
         `uvm_info("step_compare", $sformatf("Checked PC 0d%0d times", num_pc_checks), UVM_LOW);
      end
      else begin
         `uvm_error("step_compare", "PC was checked 0 times!");
      end
      if (num_gpr_checks > 0) begin
         `uvm_info("step_compare", $sformatf("Checked GPR 0d%0d times", num_gpr_checks), UVM_LOW);
      end
      else begin
         `uvm_error("step_compare", "GPR was checked 0 times!");
      end
      if (num_csr_checks > 0) begin
         `uvm_info("step_compare", $sformatf("Checked CSR 0d%0d times", num_csr_checks), UVM_LOW);
      end
      else begin
         `uvm_error("step_compare", "CSR was checked 0 times!");
      end
   endfunction // report_step_compare
   
endinterface: uvmt_cv32e40p_step_compare_if

// Interface to debug assertions and covergroups
interface uvmt_cv32e40p_debug_cov_assert_if
    import cv32e40p_pkg::*;
    (
    input  clk_i,
    input  rst_ni,

    // Core inputs
    input         fetch_enable_i, // external core fetch enable

    // External interrupt interface
    input  [31:0] irq_i,
    input         irq_ack_o,
    input  [4:0]  irq_id_o,
    input  [31:0] mie_q,

    // Instruction fetch stage
    input         if_stage_instr_rvalid_i, // Instruction word is valid
    input  [31:0] if_stage_instr_rdata_i, // Instruction word data

    // Instruction ID stage (determines executed instructions)  
    input         id_stage_instr_valid_i, // instruction word is valid
    input  [31:0] id_stage_instr_rdata_i, // Instruction word data
    input         id_stage_is_compressed,
    input  [31:0] id_stage_pc, // Program counter in decode
    input  [31:0] if_stage_pc, // Program counter in fetch
    input         is_decoding,
    input         branch_taken_ex_i,
    input         data_err_i,
    input         is_fetch_failed_i,
    input         id_valid,
    input wire ctrl_state_e  ctrl_fsm_cs,            // Controller FSM states with debug_req
    input         illegal_insn_i,
    input         illegal_insn_q, // output from controller
    input         ecall_insn_i,

    input  [31:0] boot_addr_i,

    input         rvfi_valid,
    input  [31:0] rvfi_insn,
    input         apu_req,
    input         apu_gnt,
    input         apu_busy,

    // Debug signals
    input         debug_req_i, // From controller
    input         debug_mode_q, // From controller
    input  [31:0] dcsr_q, // From controller
    input  [31:0] depc_q, // From cs regs
    input  [31:0] depc_n, // 
    input  [31:0] dm_halt_addr_i,
    input  [31:0] dm_exception_addr_i,

    input  [5:0]  mcause_q,
    input  [31:0] mtvec,
    input  [31:0] mepc_q,
    input  [31:0] tdata1,
    input  [31:0] tdata2,
    input  trigger_match_i,

    // Counter related input from cs_registers
    input  [31:0] mcountinhibit_q,
    input  [63:0] mcycle,
    input  [63:0] minstret,
    input  inst_ret,
    // WFI Interface
    input  core_sleep_o,

    input  fence_i,
      
    input  csr_access,
    input  [1:0] csr_op,
    input  [1:0] csr_op_dec,
    input  [11:0] csr_addr,
    input  csr_we_int,

    output logic is_wfi,
    output logic in_wfi,
    output logic dpc_will_hit,
    output logic addr_match,
    output logic is_ebreak,
    output logic is_cebreak,
    output logic is_dret,
    output logic is_mulhsu,
    output logic [31:0] pending_enabled_irq,
    input  pc_set,
    input  branch_in_decode
);

  clocking mon_cb @(posedge clk_i);    
    input #1step
    fetch_enable_i,

    irq_i,
    irq_ack_o,
    irq_id_o,
    mie_q,

    if_stage_instr_rvalid_i,
    if_stage_instr_rdata_i,

    id_stage_instr_valid_i,
    id_stage_instr_rdata_i,
    id_stage_is_compressed,
    id_stage_pc,
    if_stage_pc,
    is_decoding,
    branch_taken_ex_i,
    is_fetch_failed_i,
    id_valid,
    ctrl_fsm_cs,
    illegal_insn_i,
    illegal_insn_q,
    ecall_insn_i,
    boot_addr_i,
    rvfi_valid,
    rvfi_insn,
    apu_req,
    apu_gnt,
    apu_busy,
    debug_req_i,
    debug_mode_q,
    dcsr_q,
    depc_q,
    depc_n,
    dm_halt_addr_i,
    dm_exception_addr_i,
    mcause_q,
    mtvec,
    mepc_q,
    tdata1,
    tdata2,
    trigger_match_i,
    fence_i,
    mcountinhibit_q,
    mcycle,
    minstret,
    inst_ret,
    
    core_sleep_o,
    csr_access,
    csr_op,
    csr_op_dec,
    csr_addr,
    is_wfi,
    in_wfi,
    dpc_will_hit,
    addr_match,
    is_ebreak,
    is_cebreak,
    is_dret,
    is_mulhsu,
    pending_enabled_irq,
    pc_set,
    branch_in_decode;
  endclocking : mon_cb

endinterface : uvmt_cv32e40p_debug_cov_assert_if


// core-v-verif simplify rvvi for coverage collection purpose 
  `define DEF_CSR_PORTS(CSR_NAME) \
  input logic [(XLEN-1):0] csr_``CSR_NAME``_rmask, \
  input logic [(XLEN-1):0] csr_``CSR_NAME``_wmask, \
  input logic [(XLEN-1):0] csr_``CSR_NAME``_rdata, \
  input logic [(XLEN-1):0] csr_``CSR_NAME``_wdata,

  `define DEF_CSR_PORTS_VEC(CSR_NAME, VEC_SIZE) \
  input logic [(``VEC_SIZE``-1):0][(XLEN-1):0] csr_``CSR_NAME``_rmask, \
  input logic [(``VEC_SIZE``-1):0][(XLEN-1):0] csr_``CSR_NAME``_wmask, \
  input logic [(``VEC_SIZE``-1):0][(XLEN-1):0] csr_``CSR_NAME``_rdata, \
  input logic [(``VEC_SIZE``-1):0][(XLEN-1):0] csr_``CSR_NAME``_wdata,

  `define ASSIGN_CSR_N_WB(CSR_ADDR, CSR_NAME) \
    bit csr_``CSR_NAME``_wb; \
    wire [31:0] csr_``CSR_NAME``_w; \
    wire [31:0] csr_``CSR_NAME``_r; \
    assign csr_``CSR_NAME``_w = csr_``CSR_NAME``_wdata &   csr_``CSR_NAME``_wmask; \
    assign csr_``CSR_NAME``_r = csr_``CSR_NAME``_rdata & ~(csr_``CSR_NAME``_wmask); \
    assign csr[``CSR_ADDR]    = csr_``CSR_NAME``_w | csr_``CSR_NAME``_r; \
    assign csr_wb[``CSR_ADDR] = csr_``CSR_NAME``_wb; \
    always @(csr[``CSR_ADDR]) begin \
        csr_``CSR_NAME``_wb = 1; \
    end \
    always @(posedge clk) begin \
        if (valid && csr_``CSR_NAME``_wb) begin \
            csr_``CSR_NAME``_wb = 0; \
        end \
    end

  `define ASSIGN_CSR_N_WB_VEC(CSR_ADDR, CSR_NAME, CSR_ID) \
    bit csr_``CSR_NAME`` ``CSR_ID``_wb; \
    wire [31:0] csr_``CSR_NAME`` ``CSR_ID``_w; \
    wire [31:0] csr_``CSR_NAME`` ``CSR_ID``_r; \
    assign csr_``CSR_NAME`` ``CSR_ID``_w = csr_``CSR_NAME``_wdata[``CSR_ID] &   csr_``CSR_NAME``_wmask[``CSR_ID]; \
    assign csr_``CSR_NAME`` ``CSR_ID``_r = csr_``CSR_NAME``_rdata[``CSR_ID] & ~(csr_``CSR_NAME``_wmask[``CSR_ID]); \
    assign csr[``CSR_ADDR]              = csr_``CSR_NAME`` ``CSR_ID``_w | csr_``CSR_NAME`` ``CSR_ID``_r; \
    assign csr_wb[``CSR_ADDR]           = csr_``CSR_NAME`` ``CSR_ID``_wb; \
    always @(csr[``CSR_ADDR]) begin \
        csr_``CSR_NAME`` ``CSR_ID``_wb = 1; \
    end \
    always @(posedge clk) begin \
        if (valid && csr_``CSR_NAME`` ``CSR_ID``_wb) begin \
            csr_``CSR_NAME`` ``CSR_ID``_wb = 0; \
        end \
    end

interface uvmt_cv32e40p_rvvi_if #(
  parameter int ILEN    = 32,
  parameter int XLEN    = 32
) (
    
  input                               clk,
  input                               valid,
  input logic [(ILEN-1):0]            insn,
  input                               trap,
  input logic [31:0]                  pc_rdata,
  input logic [31:0]                  wa_csr_mip,

  uvma_interrupt_if                   interrupt_if,
  uvma_debug_if                       debug_if,

  // Currently only define specific csrs for current usage
  `DEF_CSR_PORTS(lpstart0)
  `DEF_CSR_PORTS(lpend0)
  `DEF_CSR_PORTS(lpcount0)
  `DEF_CSR_PORTS(lpstart1)
  `DEF_CSR_PORTS(lpend1)
  `DEF_CSR_PORTS(lpcount1)
  `DEF_CSR_PORTS(mstatus)
  `DEF_CSR_PORTS(mie)
  `DEF_CSR_PORTS(mtvec)
  `DEF_CSR_PORTS(mcause)
  `DEF_CSR_PORTS(mip)
  `DEF_CSR_PORTS(dcsr)
  `DEF_CSR_PORTS_VEC(tdata,4)

  input logic [31:0]                  dm_halt_addr
 
);

  wire [31:0]                 valid_irq;
  wire [4095:0][32:0]         csr;
  wire [4095:0]               csr_wb;
  wire [4:0]                  csr_mcause_ecp_code;
  wire [2:0]                  csr_dcsr_cause;
  wire [31:0]                 csr_trig_pc;

  logic [31:0]                irq_onehot_priority;
  logic [31:0]                mtvec_base_addr;
  logic [31:0]                mip;

  // assign valid_irq            = csr[`CSR_MIP_ADDR] & csr[`CSR_MIE_ADDR]; // fixme: rvfi misses mip (pending rvfi fixes; workaround probe rtl signals - wa_csr_mip)
  assign valid_irq            = wa_csr_mip & csr[`CSR_MIE_ADDR];
  assign dbg_req              = debug_if.debug_req;
  assign mie                  = csr[`CSR_MSTATUS_ADDR][3];
  assign mip                  = csr[`CSR_MIP_ADDR];

  assign csr_mcause_irq       = csr[`CSR_MCAUSE_ADDR][31];
  assign csr_mcause_ecp_code  = csr[`CSR_MCAUSE_ADDR][4:0];
  assign csr_dcsr_ebreakm     = csr[`CSR_DCSR_ADDR][15];
  assign csr_dcsr_stepie      = csr[`CSR_DCSR_ADDR][11];
  assign csr_dcsr_cause       = csr[`CSR_DCSR_ADDR][8:6];
  assign csr_dcsr_step        = csr[`CSR_DCSR_ADDR][2];
  assign csr_trig_execute     = csr[`CSR_TDATA1_ADDR][2];
  assign csr_trig_pc          = csr[`CSR_TDATA2_ADDR];

  assign mtvec_base_addr      = {csr[`CSR_MTVEC_ADDR][31:8], 8'h0};

  // can be expanded. Currently only define for current usage
  `ASSIGN_CSR_N_WB(`CSR_LPSTART0_ADDR, lpstart0)
  `ASSIGN_CSR_N_WB(`CSR_LPEND0_ADDR, lpend0)
  `ASSIGN_CSR_N_WB(`CSR_LPCOUNT0_ADDR, lpcount0)
  `ASSIGN_CSR_N_WB(`CSR_LPSTART1_ADDR, lpstart1)
  `ASSIGN_CSR_N_WB(`CSR_LPEND1_ADDR, lpend1)
  `ASSIGN_CSR_N_WB(`CSR_LPCOUNT1_ADDR, lpcount1)
  `ASSIGN_CSR_N_WB(`CSR_MSTATUS_ADDR, mstatus)
  `ASSIGN_CSR_N_WB(`CSR_MIE_ADDR, mie)
  `ASSIGN_CSR_N_WB(`CSR_MTVEC_ADDR, mtvec)
  `ASSIGN_CSR_N_WB(`CSR_MCAUSE_ADDR, mcause)
  `ASSIGN_CSR_N_WB(`CSR_MIP_ADDR, mip)
  `ASSIGN_CSR_N_WB(`CSR_DCSR_ADDR, dcsr)
  //`ASSIGN_CSR_N_WB_VEC(`CSR_TDATA1_ADDR, tdata, 1);
  //`ASSIGN_CSR_N_WB_VEC(`CSR_TDATA2_ADDR, tdata, 2);

  // irq_onehot_priority assignment (refer cv32e40p user manual, section 10.2)
  // priority order (high->low) is irq[31]...irq[16], irq[11], irq[3], irq[7]
  always @(valid_irq) begin
    irq_onehot_priority = 0;
    for (int i = 31; i != 0; i--) begin
      if (valid_irq[i] && (i inside {31,30,29,28,27,26,25,24,23,22,21,20,19,18,17,16, 11,3,7})) begin
        if (i == 7 && valid_irq[3]) continue;
        else begin irq_onehot_priority[i] = valid_irq[i]; break; end
      end
    end
  end
    
endinterface

//
//Interface for custom TB coverage component
//
interface uvmt_cv32e40p_cov_if

  import uvm_pkg::*;
  import uvme_cv32e40p_pkg::*;
  (
    input               clk_i,
    input               rst_ni,
    input               if_stage_instr_rvalid_i,
    input  [31:0]       if_stage_instr_rdata_i,
    input               id_stage_instr_valid_i,
    input               id_stage_id_valid_o,
    input  [31:0]       id_stage_instr_rdata_i,
    input               apu_req,
    input               apu_gnt,
    input               apu_busy,
    input  [5:0]        apu_op,
    input               apu_rvalid_i,
    input               apu_perf_wb_o,
    input  [5:0]        id_stage_apu_op_ex_o,
    input               id_stage_apu_en_ex_o,
    input  [5:0]        regfile_waddr_wb_o,  // regfile write port A addr from WB stage (lsu write-back)
    input               regfile_we_wb_o,
    input  [5:0]        regfile_alu_waddr_ex_o, // regfile write port B addr from EX stage (forwarding)
    input               regfile_alu_we_ex_o,
    input               ex_mulh_active,
    input  [2:0]        ex_mult_op_ex,
    input               ex_data_misaligned_i,
    input               ex_data_misaligned_ex_i,
    input               ex_data_req_i,
    input               ex_data_rvalid_i,
    input               ex_regfile_alu_we_i,
    input               ex_apu_valid,
    input               ex_apu_rvalid_q,
    input               debug_req_i,
    input               debug_mode_q,
    input  [31:0]       dcsr_q,
    input               trigger_match_i,

    output logic[5:0]   o_curr_fpu_apu_op_if,
    output logic[5:0]   o_last_fpu_apu_op_if,
    output logic[4:0]   if_clk_cycle_window,
    output [4:0]        curr_fpu_fd,
    output [4:0]        curr_fpu_rd,
    output [5:0]        curr_rd_at_ex_regfile_wr_contention,
    output [5:0]        curr_rd_at_wb_regfile_wr_contention,
    output [5:0]        prev_rd_waddr_contention,
    output logic[1:0]   contention_state,
    output              b2b_contention,
    output              is_mulh_ex,
    output              is_misaligned_data_req_ex,
    output              is_post_inc_ld_st_inst_ex,
    output              ex_apu_valid_memorised
  );

  `ifdef FPU_ADDMUL_LAT
  parameter int FPU_LAT_1_CYC = `FPU_ADDMUL_LAT;
  `else
  parameter int FPU_LAT_1_CYC = 0;
  `endif

  logic [4:0]       clk_cycle_window;
  logic [5:0]       curr_fpu_apu_op_if;
  logic [5:0]       last_fpu_contention_op_if;
  logic [5:0]       prev_regfile_waddr_contention;
  logic [4:0]       regfile_waddr_wb_fd;
  logic [4:0]       regfile_alu_waddr_ex_fd;
  logic [4:0]       regfile_waddr_wb_rd;
  logic [4:0]       regfile_alu_waddr_ex_rd;
  logic [5:0]       regfile_waddr_ex_contention;
  logic [5:0]       regfile_waddr_wb_contention;
  logic [1:0]       contention_valid;
  logic             b2b_contention_valid;
  logic [31:0]      current_instr_rdata;
  logic [31:0]      previous_instr_rdata;

  initial begin
      clk_cycle_window = 0;
      curr_fpu_apu_op_if = 0;
      regfile_waddr_wb_fd = 0;
      regfile_alu_waddr_ex_fd = 0;
      regfile_waddr_wb_rd = 0;
      regfile_alu_waddr_ex_rd = 0;
      regfile_waddr_ex_contention = 0;
      regfile_waddr_wb_contention = 0;
      contention_valid = 0;
      b2b_contention_valid = 0;
  end

  clocking mon_cb @(posedge clk_i);
      default input #1step output #1ns;
      input if_stage_instr_rvalid_i;
      input if_stage_instr_rdata_i;
      input id_stage_instr_valid_i;
      input id_stage_id_valid_o;
      input id_stage_instr_rdata_i;
      input apu_req;
      input apu_gnt;
      input apu_busy;
      input apu_op;
      input apu_rvalid_i;
      input apu_perf_wb_o;
      input id_stage_apu_op_ex_o;
      input id_stage_apu_en_ex_o;
      input debug_req_i;
      input debug_mode_q;
      input trigger_match_i;
      input dcsr_q;
      inout is_mulh_ex;
      inout is_misaligned_data_req_ex;
      inout is_post_inc_ld_st_inst_ex;
      inout ex_apu_valid_memorised;
  endclocking : mon_cb

  // bhv_logic_1
  // calculate each APU operation's current clock cycle number during execution for functional coverage use
  // input(s): apu_op, 
  always @(posedge clk_i or negedge rst_ni) begin
      if(!rst_ni) begin
          clk_cycle_window = 0;
          curr_fpu_apu_op_if = 0;
      end
      else begin
          if((clk_cycle_window == 0) && (apu_req == 1)) begin
              clk_cycle_window = 1;
              curr_fpu_apu_op_if = apu_op;
          end
          else if((clk_cycle_window != 0) && (apu_req == 1)) begin
              clk_cycle_window = 1;
              curr_fpu_apu_op_if = apu_op;
          end
          else if((clk_cycle_window != 0) && (apu_busy == 1)) begin
              clk_cycle_window += 1;
          end
          else begin
              clk_cycle_window = 0;
          end
      end
  end

  // bhv_logic_1a
  // sample decoded instr that execute in progress
  always @(posedge clk_i or negedge rst_ni) begin
    if(!rst_ni) begin
      previous_instr_rdata <= 0;
      current_instr_rdata  <= 0;
    end
    else begin
      if (id_stage_instr_valid_i && id_stage_id_valid_o) begin
        previous_instr_rdata <= current_instr_rdata;
        current_instr_rdata  <= id_stage_instr_rdata_i;
      end
      else begin
        previous_instr_rdata <= current_instr_rdata;
      end
    end
  end

  // bhv_logic_2 (revised)
  // Model APU contention state in EX/WB for functional coverage
  // input(s): apu_perf_wb_o, regfile_waddr_wb_o, regfile_alu_waddr_ex_o
  always @(posedge clk_i or negedge rst_ni) begin
      if(!rst_ni) begin
          contention_valid <= 0;
          b2b_contention_valid <= 0;
          last_fpu_contention_op_if <= 0;
          prev_regfile_waddr_contention <= 0;
      end
      else begin
          if (((contention_valid == 0) || (contention_valid == 2)) && (apu_perf_wb_o)) begin
            contention_valid <= 1; //set contention_valid
            b2b_contention_valid <= 0;
            last_fpu_contention_op_if <= curr_fpu_apu_op_if;
          end
          else if((contention_valid == 1) && (apu_perf_wb_o)) begin
            contention_valid <= 1; //reset contention_valid
            b2b_contention_valid <= 1;
            // if no APU execution during contention then nothing to do
            // during contention another APU transaction cannot go through
          end
          else if((contention_valid == 1) && (!apu_perf_wb_o)) begin
              contention_valid <= 2; //stalled write complete after contention
              b2b_contention_valid <= 1;
              if (FPU_LAT_1_CYC != 1) begin // IS_0_OR_2_CYCLAT
                prev_regfile_waddr_contention <= regfile_alu_waddr_ex_o; // port B
              end
              else begin // IS_1_CYCLAT
                prev_regfile_waddr_contention <= regfile_waddr_wb_o; // port A
              end
          end
          else begin
              contention_valid <= 0;
              b2b_contention_valid <= 0;
              prev_regfile_waddr_contention <= 0;
          end
      end
  end


  // bhv_logic_3
  // sample each APU operation's destination register address for functional coverage
  // input(s): apu_req, apu_busy, regfile_alu_we_ex_o, regfile_we_wb_o,  apu_rvalid_i
  always @(posedge clk_i or negedge rst_ni) begin
      if(!rst_ni) begin
          regfile_alu_waddr_ex_fd <= 0;
          regfile_alu_waddr_ex_rd <= 0;
          regfile_waddr_wb_fd <= 0;
          regfile_waddr_wb_rd <= 0;
          regfile_waddr_wb_contention <= 0;
          regfile_waddr_ex_contention <= 0;
      end
      else begin
        if (FPU_LAT_1_CYC != 1) begin // IS_0_OR_2_CYCLAT
          //Case for FPU Latency {0,2,3,4}, with regfile write from EX stage with highest priority of APU
          if (((apu_req == 1) || (apu_busy == 1)) && (regfile_alu_we_ex_o == 1) && (apu_rvalid_i == 1)) begin
              regfile_alu_waddr_ex_fd <= (regfile_alu_waddr_ex_o - 32);
              regfile_alu_waddr_ex_rd <= (regfile_alu_waddr_ex_o < 32) ? regfile_alu_waddr_ex_o : 0;
              regfile_waddr_ex_contention <= 0;
              regfile_waddr_wb_contention <= 0;
          end
          else if ((contention_valid == 1) && (regfile_alu_we_ex_o == 1) && !apu_perf_wb_o) begin // write for stalled regfile wr at contention
              regfile_alu_waddr_ex_fd <= 0;
              regfile_alu_waddr_ex_rd <= 0;
              regfile_waddr_ex_contention <= regfile_alu_waddr_ex_o; //should not be >31, check for illegal in coverage
              regfile_waddr_wb_contention <= 0;
          end
          else begin
              regfile_alu_waddr_ex_fd <= 0;
              regfile_alu_waddr_ex_rd <= 0;
              regfile_waddr_wb_fd <= 0;
              regfile_waddr_wb_rd <= 0;
              regfile_waddr_ex_contention <= 0;
              regfile_waddr_wb_contention <= 0;
          end
        end // IS_0_OR_2_CYCLAT
        else begin // IS_1_CYCLAT
          //Case FPU Latency = 1; regfile wr from WB;LSU > priority;no LSU contention, F-inst regfile wr succeed
          if ((apu_busy == 1) && (regfile_we_wb_o == 1) && (apu_rvalid_i == 1) && (!apu_perf_wb_o)) begin
              regfile_waddr_wb_fd <= (regfile_waddr_wb_o - 32);
              regfile_waddr_wb_rd <= (regfile_waddr_wb_o < 32) ? regfile_waddr_wb_o : 0;
              regfile_waddr_ex_contention <= 0;
              regfile_waddr_wb_contention <= 0;
          end
          //Case FPU Latency = 1; regfile wr from WB;LSU > priority;LSU contention,F-inst regfile wr stall
          else if((apu_busy == 1) && (regfile_we_wb_o == 1) && (apu_rvalid_i == 1) && (apu_perf_wb_o)) begin
              regfile_waddr_wb_fd <= 0;
              regfile_waddr_wb_rd <= 0;
              regfile_waddr_ex_contention <= 0;
              regfile_waddr_wb_contention = regfile_waddr_wb_o; //should not be >31, check for illegal in coverage
          end
          //Case FPU Latency = 1;regfile wr from WB;LSU > priority;LSU contention - FPU reg write cycle after contention
          else if((contention_valid == 1) && (regfile_we_wb_o == 1) && !apu_perf_wb_o) begin
              regfile_waddr_wb_fd <= (regfile_waddr_wb_o - 32);
              regfile_waddr_wb_rd <= (regfile_waddr_wb_o < 32) ? regfile_waddr_wb_o : 0;
              regfile_waddr_ex_contention <= 0;
              regfile_waddr_wb_contention <= 0;
          end
          else begin
              regfile_alu_waddr_ex_fd <= 0;
              regfile_alu_waddr_ex_rd <= 0;
              regfile_waddr_wb_fd <= 0;
              regfile_waddr_wb_rd <= 0;
              regfile_waddr_ex_contention <= 0;
              regfile_waddr_wb_contention <= 0;
          end
        end // IS_1_CYCLAT
      end
  end

  assign curr_fpu_fd = regfile_alu_waddr_ex_fd | regfile_waddr_wb_fd;
  assign curr_fpu_rd = regfile_alu_waddr_ex_rd | regfile_waddr_wb_rd;
  assign if_clk_cycle_window = clk_cycle_window;
  assign o_curr_fpu_apu_op_if = curr_fpu_apu_op_if;
  assign o_last_fpu_apu_op_if = last_fpu_contention_op_if;
  assign curr_rd_at_ex_regfile_wr_contention = regfile_waddr_ex_contention;
  assign curr_rd_at_wb_regfile_wr_contention = regfile_waddr_wb_contention;
  assign contention_state = contention_valid;
  assign b2b_contention = b2b_contention_valid;
  assign prev_rd_waddr_contention = prev_regfile_waddr_contention;
  assign is_mulh_ex = ex_mulh_active && (ex_mult_op_ex == 3'h6);
  assign is_misaligned_data_req_ex = ex_data_misaligned_i || ex_data_misaligned_ex_i;
  assign is_post_inc_ld_st_inst_ex = (ex_data_req_i || ex_data_rvalid_i) && ex_regfile_alu_we_i;
  assign ex_apu_valid_memorised = ex_apu_valid & ex_apu_rvalid_q;

endinterface : uvmt_cv32e40p_cov_if

`endif // __UVMT_CV32E40P_TB_IFS_SV__
