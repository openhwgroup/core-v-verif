`define  FORMAL  1
