//
// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2020 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//


`ifndef __UVMT_CV32E40S_TB_SV__
`define __UVMT_CV32E40S_TB_SV__


/**
 * Module encapsulating the CV32E40S DUT wrapper, and associated SV interfaces.
 * Also provide UVM environment entry and exit points.
 */
`default_nettype none
module uvmt_cv32e40s_tb;

   import uvm_pkg::*;
   import cv32e40s_pkg::*;
   import uvmt_cv32e40s_pkg::*;
   import uvme_cv32e40s_pkg::*;

   // ENV (testbench) parameters
   parameter int ENV_PARAM_INSTR_ADDR_WIDTH  = 32;
   parameter int ENV_PARAM_INSTR_DATA_WIDTH  = 32;
   parameter int ENV_PARAM_RAM_ADDR_WIDTH    = 22;

   // Capture regs for test status from Virtual Peripheral in dut_wrap.mem_i
   bit        tp;
   bit        tf;
   bit        evalid;
   bit [31:0] evalue;

   // Agent interfaces
   uvma_isacov_if               isacov_if();
   uvma_clknrst_if              clknrst_if(); // clock and resets from the clknrst agent
   uvma_clknrst_if              clknrst_if_iss();
   uvma_debug_if                debug_if();
   uvma_interrupt_if            interrupt_if();
   uvma_clic_if                 clic_if();
   uvma_obi_memory_if           obi_instr_if_i(
     .clk(clknrst_if.clk),
     .reset_n(clknrst_if.reset_n)
   );
   uvma_obi_memory_if           obi_data_if_i(
     .clk(clknrst_if.clk),
     .reset_n(clknrst_if.reset_n)
   );
   uvma_fencei_if               fencei_if_i(
     .clk(clknrst_if.clk),
     .reset_n(clknrst_if.reset_n)
   );

   // DUT Wrapper Interfaces
   uvmt_cv32e40s_vp_status_if       vp_status_if(.tests_passed(),
                                                 .tests_failed(),
                                                 .exit_valid(),
                                                 .exit_value()); // Status information generated by the Virtual Peripherals in the DUT WRAPPER memory.
   uvme_cv32e40s_core_cntrl_if      core_cntrl_if();
   uvmt_cv32e40s_core_status_if     core_status_if(.core_busy(),
                                                   .sec_lvl());     // Core status outputs

  /**
   * DUT WRAPPER instance:
   * This is an update of the riscv_wrapper.sv from PULP-Platform RI5CY project with
   * a few mods to bring unused ports from the CORE to this level using SV interfaces.
   */
   uvmt_cv32e40s_dut_wrap  #(
                             .B_EXT             (uvmt_cv32e40s_pkg::B_EXT),
                             .PMA_NUM_REGIONS   (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_NUM_REGIONS),
                             .PMA_CFG           (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_CFG),
                             .PMP_GRANULARITY   (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_GRANULARITY),
                             .PMP_NUM_REGIONS   (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_NUM_REGIONS),
                             .INSTR_ADDR_WIDTH  (ENV_PARAM_INSTR_ADDR_WIDTH),
                             .INSTR_RDATA_WIDTH (ENV_PARAM_INSTR_DATA_WIDTH),
                             .RAM_ADDR_WIDTH    (ENV_PARAM_RAM_ADDR_WIDTH),
                             .SMCLIC            (uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC)
                            )
                            dut_wrap (
                              .clknrst_if(clknrst_if),
                              .interrupt_if(interrupt_if),
                              .vp_status_if(vp_status_if),
                              .core_cntrl_if(core_cntrl_if),
                              .core_status_if(core_status_if),
                              .obi_instr_if_i(obi_instr_if_i),
                              .obi_data_if_i(obi_data_if_i),
                              .fencei_if_i(fencei_if_i),
                              .clic_if(clic_if),
                              .*);

  bind cv32e40s_wrapper
    uvma_rvfi_instr_if#(uvme_cv32e40s_pkg::ILEN,
                        uvme_cv32e40s_pkg::XLEN) rvfi_instr_if_0_i(.clk(clk_i),
                                                                   .reset_n(rst_ni),

                                                                   .rvfi_valid(rvfi_i.rvfi_valid[0]),
                                                                   .rvfi_order(rvfi_i.rvfi_order[uvma_rvfi_pkg::ORDER_WL*0+:uvma_rvfi_pkg::ORDER_WL]),
                                                                   .rvfi_insn(rvfi_i.rvfi_insn[uvme_cv32e40s_pkg::ILEN*0+:uvme_cv32e40s_pkg::ILEN]),
                                                                   .rvfi_trap(rvfi_i.rvfi_trap[11:0]),
                                                                   .rvfi_halt(rvfi_i.rvfi_halt[0]),
                                                                   .rvfi_intr(rvfi_i.rvfi_intr),
                                                                   .rvfi_dbg(rvfi_i.rvfi_dbg),
                                                                   .rvfi_dbg_mode(rvfi_i.rvfi_dbg_mode),
                                                                   .rvfi_nmip(rvfi_i.rvfi_nmip),
                                                                   .rvfi_mode(rvfi_i.rvfi_mode[uvma_rvfi_pkg::MODE_WL*0+:uvma_rvfi_pkg::MODE_WL]),
                                                                   .rvfi_ixl(rvfi_i.rvfi_ixl[uvma_rvfi_pkg::IXL_WL*0+:uvma_rvfi_pkg::IXL_WL]),
                                                                   .rvfi_pc_rdata(rvfi_i.rvfi_pc_rdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_pc_wdata(rvfi_i.rvfi_pc_wdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rs1_addr(rvfi_i.rvfi_rs1_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
                                                                   .rvfi_rs1_rdata(rvfi_i.rvfi_rs1_rdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rs2_addr(rvfi_i.rvfi_rs2_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
                                                                   .rvfi_rs2_rdata(rvfi_i.rvfi_rs2_rdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rs3_addr('0),
                                                                   .rvfi_rs3_rdata('0),
                                                                   .rvfi_rd1_addr(rvfi_i.rvfi_rd_addr[uvma_rvfi_pkg::GPR_ADDR_WL*0+:uvma_rvfi_pkg::GPR_ADDR_WL]),
                                                                   .rvfi_rd1_wdata(rvfi_i.rvfi_rd_wdata[uvme_cv32e40s_pkg::XLEN*0+:uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_rd2_addr('0),
                                                                   .rvfi_rd2_wdata('0),
                                                                   .rvfi_gpr_rdata(rvfi_i.rvfi_gpr_rdata[32*uvme_cv32e40s_pkg::XLEN*0  +:32*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_gpr_rmask(rvfi_i.rvfi_gpr_rmask[32*0  +:32]),
                                                                   .rvfi_gpr_wdata(rvfi_i.rvfi_gpr_wdata[32*uvme_cv32e40s_pkg::XLEN*0  +:32*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_gpr_wmask(rvfi_i.rvfi_gpr_wmask[32*0  +:32]),
                                                                   .rvfi_mem_addr(rvfi_i.rvfi_mem_addr[  uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_mem_rdata(rvfi_i.rvfi_mem_rdata[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_mem_rmask(rvfi_i.rvfi_mem_rmask[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8*0  +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8]),
                                                                   .rvfi_mem_wdata(rvfi_i.rvfi_mem_wdata[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN*0    +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN]),
                                                                   .rvfi_mem_wmask(rvfi_i.rvfi_mem_wmask[uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8*0  +:uvma_rvfi_pkg::NMEM*uvme_cv32e40s_pkg::XLEN/8])
                                                                   );

  // RVFI CSR binds
  `RVFI_CSR_BIND(marchid)
  `RVFI_CSR_BIND(mcountinhibit)
  `RVFI_CSR_BIND(mstatus)
  `RVFI_CSR_BIND(mstatush)
  `RVFI_CSR_BIND(mcounteren)
  `RVFI_CSR_BIND(menvcfg)
  `RVFI_CSR_BIND(menvcfgh)
  `RVFI_CSR_BIND(mvendorid)
  `RVFI_CSR_BIND(misa)
  `RVFI_CSR_BIND(mtvec)
  `RVFI_CSR_BIND(mtval)
  `RVFI_CSR_BIND(mscratch)
  `RVFI_CSR_BIND(mepc)
  `RVFI_CSR_BIND(mcause)
  `RVFI_CSR_BIND(mip)
  `RVFI_CSR_BIND(mie)
  `RVFI_CSR_BIND(mhartid)
  `RVFI_CSR_BIND(mimpid)
  `RVFI_CSR_BIND(minstret)
  `RVFI_CSR_BIND(minstreth)
  `RVFI_CSR_BIND(mcycle)
  `RVFI_CSR_BIND(mcycleh)

  `RVFI_CSR_BIND(dcsr)
  `RVFI_CSR_BIND(dpc)
  `RVFI_CSR_BIND(tselect)
  `RVFI_CSR_BIND(tinfo)

  `RVFI_CSR_IDX_BIND(mhpmcounter,,3)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,4)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,5)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,6)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,7)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,8)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,9)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,10)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,11)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,12)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,13)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,14)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,15)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,16)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,17)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,18)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,19)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,20)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,21)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,22)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,23)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,24)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,25)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,26)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,27)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,28)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,29)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,30)
  `RVFI_CSR_IDX_BIND(mhpmcounter,,31)

  `RVFI_CSR_IDX_BIND(pmpcfg,,0)
  `RVFI_CSR_IDX_BIND(pmpcfg,,1)
  `RVFI_CSR_IDX_BIND(pmpcfg,,2)
  `RVFI_CSR_IDX_BIND(pmpcfg,,3)
  `RVFI_CSR_IDX_BIND(pmpcfg,,4)
  `RVFI_CSR_IDX_BIND(pmpcfg,,5)
  `RVFI_CSR_IDX_BIND(pmpcfg,,6)
  `RVFI_CSR_IDX_BIND(pmpcfg,,7)
  `RVFI_CSR_IDX_BIND(pmpcfg,,8)
  `RVFI_CSR_IDX_BIND(pmpcfg,,9)
  `RVFI_CSR_IDX_BIND(pmpcfg,,10)
  `RVFI_CSR_IDX_BIND(pmpcfg,,11)
  `RVFI_CSR_IDX_BIND(pmpcfg,,12)
  `RVFI_CSR_IDX_BIND(pmpcfg,,13)
  `RVFI_CSR_IDX_BIND(pmpcfg,,14)
  `RVFI_CSR_IDX_BIND(pmpcfg,,15)

  `RVFI_CSR_IDX_BIND(pmpaddr,,0)
  `RVFI_CSR_IDX_BIND(pmpaddr,,1)
  `RVFI_CSR_IDX_BIND(pmpaddr,,2)
  `RVFI_CSR_IDX_BIND(pmpaddr,,3)
  `RVFI_CSR_IDX_BIND(pmpaddr,,4)
  `RVFI_CSR_IDX_BIND(pmpaddr,,5)
  `RVFI_CSR_IDX_BIND(pmpaddr,,6)
  `RVFI_CSR_IDX_BIND(pmpaddr,,7)
  `RVFI_CSR_IDX_BIND(pmpaddr,,8)
  `RVFI_CSR_IDX_BIND(pmpaddr,,9)
  `RVFI_CSR_IDX_BIND(pmpaddr,,10)
  `RVFI_CSR_IDX_BIND(pmpaddr,,11)
  `RVFI_CSR_IDX_BIND(pmpaddr,,12)
  `RVFI_CSR_IDX_BIND(pmpaddr,,13)
  `RVFI_CSR_IDX_BIND(pmpaddr,,14)
  `RVFI_CSR_IDX_BIND(pmpaddr,,15)
  `RVFI_CSR_IDX_BIND(pmpaddr,,16)
  `RVFI_CSR_IDX_BIND(pmpaddr,,17)
  `RVFI_CSR_IDX_BIND(pmpaddr,,18)
  `RVFI_CSR_IDX_BIND(pmpaddr,,19)
  `RVFI_CSR_IDX_BIND(pmpaddr,,20)
  `RVFI_CSR_IDX_BIND(pmpaddr,,21)
  `RVFI_CSR_IDX_BIND(pmpaddr,,22)
  `RVFI_CSR_IDX_BIND(pmpaddr,,23)
  `RVFI_CSR_IDX_BIND(pmpaddr,,24)
  `RVFI_CSR_IDX_BIND(pmpaddr,,25)
  `RVFI_CSR_IDX_BIND(pmpaddr,,26)
  `RVFI_CSR_IDX_BIND(pmpaddr,,27)
  `RVFI_CSR_IDX_BIND(pmpaddr,,28)
  `RVFI_CSR_IDX_BIND(pmpaddr,,29)
  `RVFI_CSR_IDX_BIND(pmpaddr,,30)
  `RVFI_CSR_IDX_BIND(pmpaddr,,31)
  `RVFI_CSR_IDX_BIND(pmpaddr,,32)
  `RVFI_CSR_IDX_BIND(pmpaddr,,33)
  `RVFI_CSR_IDX_BIND(pmpaddr,,34)
  `RVFI_CSR_IDX_BIND(pmpaddr,,35)
  `RVFI_CSR_IDX_BIND(pmpaddr,,36)
  `RVFI_CSR_IDX_BIND(pmpaddr,,37)
  `RVFI_CSR_IDX_BIND(pmpaddr,,38)
  `RVFI_CSR_IDX_BIND(pmpaddr,,39)
  `RVFI_CSR_IDX_BIND(pmpaddr,,40)
  `RVFI_CSR_IDX_BIND(pmpaddr,,41)
  `RVFI_CSR_IDX_BIND(pmpaddr,,42)
  `RVFI_CSR_IDX_BIND(pmpaddr,,43)
  `RVFI_CSR_IDX_BIND(pmpaddr,,44)
  `RVFI_CSR_IDX_BIND(pmpaddr,,45)
  `RVFI_CSR_IDX_BIND(pmpaddr,,46)
  `RVFI_CSR_IDX_BIND(pmpaddr,,47)
  `RVFI_CSR_IDX_BIND(pmpaddr,,48)
  `RVFI_CSR_IDX_BIND(pmpaddr,,49)
  `RVFI_CSR_IDX_BIND(pmpaddr,,50)
  `RVFI_CSR_IDX_BIND(pmpaddr,,51)
  `RVFI_CSR_IDX_BIND(pmpaddr,,52)
  `RVFI_CSR_IDX_BIND(pmpaddr,,53)
  `RVFI_CSR_IDX_BIND(pmpaddr,,54)
  `RVFI_CSR_IDX_BIND(pmpaddr,,55)
  `RVFI_CSR_IDX_BIND(pmpaddr,,56)
  `RVFI_CSR_IDX_BIND(pmpaddr,,57)
  `RVFI_CSR_IDX_BIND(pmpaddr,,58)
  `RVFI_CSR_IDX_BIND(pmpaddr,,59)
  `RVFI_CSR_IDX_BIND(pmpaddr,,60)
  `RVFI_CSR_IDX_BIND(pmpaddr,,61)
  `RVFI_CSR_IDX_BIND(pmpaddr,,62)
  `RVFI_CSR_IDX_BIND(pmpaddr,,63)

  `RVFI_CSR_IDX_BIND(mhpmevent,,3)
  `RVFI_CSR_IDX_BIND(mhpmevent,,4)
  `RVFI_CSR_IDX_BIND(mhpmevent,,5)
  `RVFI_CSR_IDX_BIND(mhpmevent,,6)
  `RVFI_CSR_IDX_BIND(mhpmevent,,7)
  `RVFI_CSR_IDX_BIND(mhpmevent,,8)
  `RVFI_CSR_IDX_BIND(mhpmevent,,9)
  `RVFI_CSR_IDX_BIND(mhpmevent,,10)
  `RVFI_CSR_IDX_BIND(mhpmevent,,11)
  `RVFI_CSR_IDX_BIND(mhpmevent,,12)
  `RVFI_CSR_IDX_BIND(mhpmevent,,13)
  `RVFI_CSR_IDX_BIND(mhpmevent,,14)
  `RVFI_CSR_IDX_BIND(mhpmevent,,15)
  `RVFI_CSR_IDX_BIND(mhpmevent,,16)
  `RVFI_CSR_IDX_BIND(mhpmevent,,17)
  `RVFI_CSR_IDX_BIND(mhpmevent,,18)
  `RVFI_CSR_IDX_BIND(mhpmevent,,19)
  `RVFI_CSR_IDX_BIND(mhpmevent,,20)
  `RVFI_CSR_IDX_BIND(mhpmevent,,21)
  `RVFI_CSR_IDX_BIND(mhpmevent,,22)
  `RVFI_CSR_IDX_BIND(mhpmevent,,23)
  `RVFI_CSR_IDX_BIND(mhpmevent,,24)
  `RVFI_CSR_IDX_BIND(mhpmevent,,25)
  `RVFI_CSR_IDX_BIND(mhpmevent,,26)
  `RVFI_CSR_IDX_BIND(mhpmevent,,27)
  `RVFI_CSR_IDX_BIND(mhpmevent,,28)
  `RVFI_CSR_IDX_BIND(mhpmevent,,29)
  `RVFI_CSR_IDX_BIND(mhpmevent,,30)
  `RVFI_CSR_IDX_BIND(mhpmevent,,31)

  `RVFI_CSR_IDX_BIND(mhpmcounter,h,3)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,4)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,5)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,6)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,7)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,8)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,9)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,10)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,11)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,12)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,13)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,14)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,15)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,16)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,17)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,18)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,19)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,20)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,21)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,22)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,23)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,24)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,25)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,26)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,27)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,28)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,29)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,30)
  `RVFI_CSR_IDX_BIND(mhpmcounter,h,31)

  `RVFI_CSR_BIND(mconfigptr)


  // dscratch0
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_dscratch0_if_0_i(.clk(clk_i),
                                                                         .reset_n(rst_ni),
                                                                         .rvfi_csr_rmask(rvfi_i.rvfi_csr_dscratch_rmask[0]),
                                                                         .rvfi_csr_wmask(rvfi_i.rvfi_csr_dscratch_wmask[0]),
                                                                         .rvfi_csr_rdata(rvfi_i.rvfi_csr_dscratch_rdata[0]),
                                                                         .rvfi_csr_wdata(rvfi_i.rvfi_csr_dscratch_wdata[0])
    );

  // dscratch1
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_dscratch1_if_0_i(.clk(clk_i),
                                                                         .reset_n(rst_ni),
                                                                         .rvfi_csr_rmask(rvfi_i.rvfi_csr_dscratch_rmask[1]),
                                                                         .rvfi_csr_wmask(rvfi_i.rvfi_csr_dscratch_wmask[1]),
                                                                         .rvfi_csr_rdata(rvfi_i.rvfi_csr_dscratch_rdata[1]),
                                                                         .rvfi_csr_wdata(rvfi_i.rvfi_csr_dscratch_wdata[1])
    );

  // tdata1
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_tdata1_if_0_i(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[1]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[1]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[1]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[1])
    );

  // tdata2
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_tdata2_if_0_i(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[2]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[2]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[2]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[2])
    );

  // tdata3
  bind cv32e40s_wrapper
    uvma_rvfi_csr_if#(uvme_cv32e40s_pkg::XLEN) rvfi_csr_tdata3_if_0_i(.clk(clk_i),
                                                                     .reset_n(rst_ni),
                                                                     .rvfi_csr_rmask(rvfi_i.rvfi_csr_tdata_rmask[3]),
                                                                     .rvfi_csr_wmask(rvfi_i.rvfi_csr_tdata_wmask[3]),
                                                                     .rvfi_csr_rdata(rvfi_i.rvfi_csr_tdata_rdata[3]),
                                                                     .rvfi_csr_wdata(rvfi_i.rvfi_csr_tdata_wdata[3])
    );

  bind uvmt_cv32e40s_dut_wrap
    uvma_obi_memory_assert_if_wrp#(
      .ADDR_WIDTH(32),
      .DATA_WIDTH(32),
      .AUSER_WIDTH(0),
      .WUSER_WIDTH(0),
      .RUSER_WIDTH(0),
      .ID_WIDTH(0),
      .ACHK_WIDTH(0),
      .RCHK_WIDTH(0),
      .IS_1P2(1)
    ) obi_instr_memory_assert_i(.obi(obi_instr_if_i));

  bind uvmt_cv32e40s_dut_wrap
    uvma_obi_memory_assert_if_wrp#(
      .ADDR_WIDTH(32),
      .DATA_WIDTH(32),
      .AUSER_WIDTH(0),
      .WUSER_WIDTH(0),
      .RUSER_WIDTH(0),
      .ID_WIDTH(0),
      .ACHK_WIDTH(0),
      .RCHK_WIDTH(0),
      .IS_1P2(1)
    ) obi_data_memory_assert_i(.obi(obi_data_if_i));

  // Bind in verification modules to the design
  `ifndef SMCLIC_EN
  bind cv32e40s_core
    uvmt_cv32e40s_interrupt_assert  interrupt_assert_i (
      .mcause_n     ({cs_registers_i.mcause_n.irq, cs_registers_i.mcause_n.exception_code[4:0]}),
      .mip          (cs_registers_i.mip_rdata),
      .mie_q        (cs_registers_i.mie_q),
      .mstatus_mie  (cs_registers_i.mstatus_q.mie),
      .mstatus_tw   (cs_registers_i.mstatus_q.tw),
      .mtvec_mode_q (cs_registers_i.mtvec_q.mode),

      .if_stage_instr_req_o    (if_stage_i.m_c_obi_instr_if.s_req.req),
      .if_stage_instr_rvalid_i (if_stage_i.m_c_obi_instr_if.s_rvalid.rvalid),
      .if_stage_instr_rdata_i  (if_stage_i.m_c_obi_instr_if.resp_payload.rdata),
      .alignbuf_outstanding    (if_stage_i.prefetch_unit_i.alignment_buffer_i.outstanding_cnt_q),

      .ex_stage_instr_valid (ex_stage_i.id_ex_pipe_i.instr_valid),

      .wb_stage_instr_valid_i    (wb_stage_i.ex_wb_pipe_i.instr_valid),
      .wb_stage_instr_rdata_i    (wb_stage_i.ex_wb_pipe_i.instr.bus_resp.rdata),
      .wb_stage_instr_err_i      (wb_stage_i.ex_wb_pipe_i.instr.bus_resp.err),
      .wb_stage_instr_mpu_status (wb_stage_i.ex_wb_pipe_i.instr.mpu_status),

      .branch_taken_ex (controller_i.controller_fsm_i.branch_taken_ex),
      .debug_mode_q    (controller_i.controller_fsm_i.debug_mode_q),

      .irq_ack_o (core_i.irq_ack),
      .irq_id_o  (core_i.irq_id),

      .*
    );
  `endif

  `ifdef SMCLIC_EN
  // CLIC assertions
  bind cv32e40s_core
    uvmt_cv32e40s_clic_interrupt_assert#(
      .SMCLIC(uvmt_cv32e40s_pkg::CORE_PARAM_SMCLIC)
    ) clic_assert_i(
      .dpc                 (cs_registers_i.dpc_rdata),
      .mintstatus          (cs_registers_i.mintstatus_rdata),
      .mintthresh          (cs_registers_i.mintthresh_rdata),
      .mcause              (cs_registers_i.mcause_rdata),
      .mtvec               (cs_registers_i.mtvec_rdata),
      .mtvt                (cs_registers_i.mtvt_rdata),
      .mclicbase           (cs_registers_i.mclicbase_rdata),
      .mepc                (cs_registers_i.mepc_rdata),
      .mip                 (cs_registers_i.mip_rdata),
      .mie                 (cs_registers_i.mie_rdata),
      .mnxti               (cs_registers_i.mnxti_rdata),
      .mscratch            (cs_registers_i.mscratch_rdata),
      .mscratchcsw         (cs_registers_i.mscratchcsw_rdata),
      .mscratchcswl        (cs_registers_i.mscratchcswl_rdata),
      .dcsr                (cs_registers_i.dcsr_rdata),

      .rvfi_mepc_wdata     (rvfi_i.rvfi_csr_mepc_wdata),
      .rvfi_mepc_wmask     (rvfi_i.rvfi_csr_mepc_wmask),
      .rvfi_mepc_rdata     (rvfi_i.rvfi_csr_mepc_rdata),
      .rvfi_mepc_rmask     (rvfi_i.rvfi_csr_mepc_rmask),
      .rvfi_dpc_rdata      (rvfi_i.rvfi_csr_dpc_rdata),
      .rvfi_dpc_rmask      (rvfi_i.rvfi_csr_dpc_rmask),
      .rvfi_mscratch_rdata (rvfi_i.rvfi_csr_mscratch_rdata),
      .rvfi_mscratch_rmask (rvfi_i.rvfi_csr_mscratch_rmask),
      .rvfi_mscratch_wdata (rvfi_i.rvfi_csr_mscratch_wdata),
      .rvfi_mscratch_wmask (rvfi_i.rvfi_csr_mscratch_wmask),

      .irq_i               (core_i.irq_i),
      .irq_ack             (core_i.irq_ack),
      .fetch_enable        (core_i.fetch_enable),
      .current_priv_mode   (core_i.priv_lvl),
      .mtvec_addr_i        (core_i.mtvec_addr_i),
      // External inputs
      .clic_if             (dut_wrap.clic_if),
      // Internal sampled   variants
      .irq_id              (core_i.irq_id[SMCLIC_ID_WIDTH-1:0]),
      .irq_level           (core_i.irq_level),
      .irq_priv            (core_i.irq_priv),
      .irq_shv             (core_i.irq_shv),

      .obi_instr_req       (core_i.instr_req_o),
      .obi_instr_gnt       (core_i.instr_gnt_i),
      .obi_instr_rvalid    (core_i.instr_rvalid_i),
      .obi_instr_addr      (core_i.instr_addr_o),
      .obi_instr_rdata     (core_i.instr_rdata_i),
      .obi_instr_rready    (1'b1),
      .obi_instr_err       (core_i.instr_err_i),

      .obi_data_addr       (core_i.data_addr_o),
      .obi_data_wdata      (core_i.data_wdata_o),
      .obi_data_we         (core_i.data_we_o),
      .obi_data_be         (core_i.data_be_o),
      .obi_data_req        (core_i.data_req_o),
      .obi_data_gnt        (core_i.data_gnt_i),
      .obi_data_rvalid     (core_i.data_rvalid_i),
      .obi_data_rready     (1'b1),
      .obi_data_err        (core_i.data_err_i),

      .debug_mode          (controller_i.controller_fsm_i.debug_mode_q),
      .debug_req           (core_i.debug_req_i),
      .debug_havereset     (core_i.debug_havereset_o),
      .debug_running       (core_i.debug_running_o),
      .debug_halt_addr     (dut_wrap.cv32e40s_wrapper_i.dm_halt_addr_i),
      .debug_exc_addr      (dut_wrap.cv32e40s_wrapper_i.dm_exception_addr_i),

      .rvfi_mode           (rvfi_i.rvfi_mode),
      .rvfi_insn           (rvfi_i.rvfi_insn),
      .rvfi_intr           (rvfi_i.rvfi_intr),
      .rvfi_rs1_rdata      (rvfi_i.rvfi_rs1_rdata),
      .rvfi_rs2_rdata      (rvfi_i.rvfi_rs2_rdata),
      .rvfi_rd_wdata       (rvfi_i.rvfi_rd_wdata),
      .rvfi_valid          (rvfi_i.rvfi_valid),
      .rvfi_pc_rdata       (rvfi_i.rvfi_pc_rdata),
      .rvfi_pc_wdata       (rvfi_i.rvfi_pc_wdata),
      .rvfi_trap           (rvfi_i.rvfi_trap),
      .rvfi_dbg_mode       (rvfi_i.rvfi_dbg_mode),
      .rvfi_dbg            (rvfi_i.rvfi_dbg),

      .wu_wfe              (dut_wrap.cv32e40s_wrapper_i.wu_wfe_i),
      .core_sleep_o        (core_i.core_sleep_o),
      .*
    );
  `endif

  // User-mode assertions

  bind  cv32e40s_wrapper
    uvmt_cv32e40s_umode_assert  umode_assert_i (
      .rvfi_valid    (rvfi_i.rvfi_valid),
      .rvfi_mode     (rvfi_i.rvfi_mode),
      .rvfi_order    (rvfi_i.rvfi_order),
      .rvfi_trap     (rvfi_i.rvfi_trap),
      .rvfi_intr     (rvfi_i.rvfi_intr),
      .rvfi_insn     (rvfi_i.rvfi_insn),
      .rvfi_dbg_mode (rvfi_i.rvfi_dbg_mode),
      .rvfi_dbg      (rvfi_i.rvfi_dbg),
      .rvfi_pc_rdata (rvfi_i.rvfi_pc_rdata),

      .rvfi_csr_dcsr_rdata       (rvfi_i.rvfi_csr_dcsr_rdata),
      .rvfi_csr_mcause_rdata     (rvfi_i.rvfi_csr_mcause_rdata),
      .rvfi_csr_mcause_wdata     (rvfi_i.rvfi_csr_mcause_wdata),
      .rvfi_csr_mcause_wmask     (rvfi_i.rvfi_csr_mcause_wmask),
      .rvfi_csr_mcounteren_rdata (rvfi_i.rvfi_csr_mcounteren_rdata),
      .rvfi_csr_misa_rdata       (rvfi_i.rvfi_csr_misa_rdata),
      .rvfi_csr_mscratch_rdata   (rvfi_i.rvfi_csr_mscratch_rdata),
      .rvfi_csr_mscratch_rmask   (rvfi_i.rvfi_csr_mscratch_rmask),
      .rvfi_csr_mscratch_wdata   (rvfi_i.rvfi_csr_mscratch_wdata),
      .rvfi_csr_mscratch_wmask   (rvfi_i.rvfi_csr_mscratch_wmask),
      .rvfi_csr_mstatus_rdata    (rvfi_i.rvfi_csr_mstatus_rdata),
      .rvfi_csr_mstatus_wdata    (rvfi_i.rvfi_csr_mstatus_wdata),
      .rvfi_csr_mstatus_wmask    (rvfi_i.rvfi_csr_mstatus_wmask),
      .rvfi_csr_mstateen0_rdata  (rvfi_i.rvfi_csr_mstateen0_rdata),

      .impu_valid (core_i.if_stage_i.mpu_i.core_trans_valid_i),
      .impu_addr  (core_i.if_stage_i.mpu_i.core_trans_i.addr),

      .*
    );

  // Fence.i assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_fencei_assert #(
      .PMA_NUM_REGIONS (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_NUM_REGIONS),
      .PMA_CFG         (uvmt_cv32e40s_pkg::CORE_PARAM_PMA_CFG)
    ) fencei_assert_i (
      .wb_valid           (core_i.wb_stage_i.wb_valid),
      .wb_instr_valid     (core_i.ex_wb_pipe.instr_valid),
      .wb_sys_en          (core_i.ex_wb_pipe.sys_en),
      .wb_sys_fencei_insn (core_i.ex_wb_pipe.sys_fencei_insn),
      .wb_pc              (core_i.ex_wb_pipe.pc),
      .wb_rdata           (core_i.ex_wb_pipe.instr.bus_resp.rdata),
      .wb_buffer_state    (core_i.load_store_unit_i.write_buffer_i.state),

      .rvfi_valid         (rvfi_i.rvfi_valid),
      .rvfi_intr          (rvfi_i.rvfi_intr.intr),
      .rvfi_dbg_mode      (rvfi_i.rvfi_dbg_mode),

      .*
    );

<<<<<<< 5524721d4a2e70904534b020a7b33efe96ac0c2a

||||||| merged common ancestors



=======
>>>>>>> Clic assertions and necessary infrastructure updates
  // Core integration assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_integration_assert  integration_assert_i (
      .*
    );


  // Xsecure assertion and coverage interface

  bind cv32e40s_wrapper
    uvmt_cv32e40s_xsecure_if  xsecure_if (

	    // Core signals: cpuctrl rdata registeret cannot be read by rvfi, we must therefore use core signales instead
      // Gated clock
      .core_clk_gated                                     (core_i.clk),

      // CSR
      .core_alert_minor_o                                 (alert_minor_o),

      .core_xsecure_ctrl_cpuctrl_dataindtiming	          (core_i.xsecure_ctrl.cpuctrl.dataindtiming),
      .core_xsecure_ctrl_cpuctrl_rnddummy		              (core_i.xsecure_ctrl.cpuctrl.rnddummy),

      .core_xsecure_ctrl_cpuctrl_rnddummyfreq             (core_i.xsecure_ctrl.cpuctrl[19:16]),
      .core_if_stage_gen_dummy_instr_dummy_instr_dummy_en (core_i.if_stage_i.gen_dummy_instr.dummy_instr_i.dummy_en),

      .core_cs_registers_xsecure_lfsr_lockup              (core_i.cs_registers_i.xsecure.lfsr_lockup),
      .core_controller_controller_fsm_debug_mode_q        (core_i.controller_i.controller_fsm_i.debug_mode_q),

      .core_cs_registers_mhpmcounter_mcycle               (core_i.cs_registers_i.mcycle_o),
      .core_cs_registers_mhpmcounter_minstret             (core_i.cs_registers_i.mhpmcounter_q[2]),
      .core_cs_registers_mhpmcounter_31_to_3              (core_i.cs_registers_i.mhpmcounter_q[31:3]),
      .core_cs_registers_mhpmevent_31_to_3                (core_i.cs_registers_i.mhpmevent_q[31:3]),
      .core_cs_registers_mcountinhibit_q_mcycle_inhibit   (core_i.cs_registers_i.mcountinhibit_q[0]),
      .core_cs_registers_mcountinhibit_q_minstret_inhibit (core_i.cs_registers_i.mcountinhibit_q[2]),

      .core_cs_registers_csr_en_gated                     (core_i.cs_registers_i.csr_en_gated),
      .core_cs_registers_csr_waddr                        (core_i.cs_registers_i.csr_waddr),

      .core_LFSR0_CFG_default_seed                        (core_i.LFSR0_CFG.default_seed),
      .core_LFSR1_CFG_default_seed                        (core_i.LFSR1_CFG.default_seed),
      .core_LFSR2_CFG_default_seed                        (core_i.LFSR2_CFG.default_seed),

      .core_xsecure_ctrl_lfsr0                            (core_i.xsecure_ctrl.lfsr0),
      .core_xsecure_ctrl_lfsr1                            (core_i.xsecure_ctrl.lfsr1),
      .core_xsecure_ctrl_lfsr2                            (core_i.xsecure_ctrl.lfsr2),

      .core_cs_registers_xsecure_lfsr0_seed_we            (core_i.cs_registers_i.xsecure.lfsr0_i.seed_we_i),
      .core_cs_registers_xsecure_lfsr1_seed_we            (core_i.cs_registers_i.xsecure.lfsr1_i.seed_we_i),
      .core_cs_registers_xsecure_lfsr2_seed_we            (core_i.cs_registers_i.xsecure.lfsr2_i.seed_we_i),

      // IF stage
      .core_if_stage_if_valid_o                           (core_i.if_stage_i.if_valid_o),
      .core_if_stage_id_ready_i                           (core_i.if_stage_i.id_ready_i),

      .core_if_stage_gen_dummy_instr_dummy_instr_lfsr_rs1 (core_i.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_rs1),
      .core_if_stage_gen_dummy_instr_dummy_instr_lfsr_rs2 (core_i.if_stage_i.gen_dummy_instr.dummy_instr_i.lfsr_rs2),

      .core_if_stage_instr_meta_n_dummy                   (core_i.if_stage_i.instr_meta_n.dummy),

      // IF ID pipe
      .core_if_id_pipe_instr_meta_dummy                   (core_i.if_id_pipe.instr_meta.dummy),
      .core_if_id_pipe_instr_bus_resp_rdata               (core_i.if_id_pipe.instr.bus_resp.rdata),

      // ID stage
      .core_id_stage_id_valid_o                           (core_i.id_stage_i.id_valid_o),
      .core_id_stage_ex_ready_i                           (core_i.id_stage_i.ex_ready_i),

      // ID EX pipe
      .core_id_ex_pipe_instr_meta_dummy                   (core_i.id_ex_pipe.instr_meta.dummy),
      .core_id_ex_pipe_instr_bus_resp_rdata               (core_i.id_ex_pipe.instr.bus_resp.rdata),

      // EX WB pipe
      .core_wb_stage_ex_wb_pipe_instr_meta_dummy          (core_i.wb_stage_i.ex_wb_pipe_i.instr_meta.dummy),

      // WB stage
      .core_wb_stage_wb_valid_o                           (core_i.wb_stage_i.wb_valid_o),
      .*
    );

    // Xsecure assertions

 bind cv32e40s_wrapper
    uvmt_cv32e40s_xsecure_assert #(
	.SECURE	(cv32e40s_pkg::SECURE)
    ) xsecure_assert_i 	(
    	.xsecure_if	(xsecure_if),
	    .rvfi_if	  (rvfi_instr_if_0_i)
    );

  // Debug assertion and coverage interface

  // Instantiate debug assertions

  bind cv32e40s_wrapper
    uvmt_cv32e40s_debug_cov_assert_if  debug_cov_assert_if (
      .id_valid               (core_i.id_stage_i.id_valid_o),
      .sys_fence_insn_i       (core_i.id_stage_i.decoder_i.sys_fencei_insn_o),

      .ex_stage_csr_en        (core_i.id_ex_pipe.csr_en),
      .ex_valid               (core_i.ex_stage_i.instr_valid),
      .ex_stage_instr_rdata_i (core_i.id_ex_pipe.instr.bus_resp.rdata),
      .ex_stage_pc            (core_i.id_ex_pipe.pc),

      .wb_stage_instr_rdata_i (core_i.ex_wb_pipe.instr.bus_resp.rdata),
      .wb_stage_instr_valid_i (core_i.ex_wb_pipe.instr_valid),
      .wb_stage_pc            (core_i.wb_stage_i.ex_wb_pipe_i.pc),
      .wb_err                 (core_i.ex_wb_pipe.instr.bus_resp.err),
      .wb_illegal             (core_i.ex_wb_pipe.illegal_insn),
      .wb_valid               (core_i.wb_stage_i.wb_valid_o),
      .wb_mpu_status          (core_i.ex_wb_pipe.instr.mpu_status),
      .illegal_insn_i         (core_i.ex_wb_pipe.illegal_insn),
      .sys_en_i               (core_i.ex_wb_pipe.sys_en),
      .sys_ecall_insn_i       (core_i.ex_wb_pipe.sys_ecall_insn),

      .ctrl_fsm_cs            (core_i.controller_i.controller_fsm_i.ctrl_fsm_cs),
      .debug_req_i            (core_i.controller_i.controller_fsm_i.debug_req_i),
      .debug_havereset        (core_i.debug_havereset_o),
      .debug_running          (core_i.debug_running_o),
      .debug_halted           (core_i.debug_halted_o),

      .debug_req_q            (core_i.controller_i.controller_fsm_i.debug_req_q),
      .pending_debug          (core_i.controller_i.controller_fsm_i.pending_debug),
      .pending_nmi            (core_i.controller_i.controller_fsm_i.pending_nmi),
      .nmi_allowed            (core_i.controller_i.controller_fsm_i.nmi_allowed),
      .debug_mode_q           (core_i.controller_i.controller_fsm_i.debug_mode_q),
      .trigger_match_in_wb    (core_i.controller_i.controller_fsm_i.trigger_match_in_wb),
      .branch_in_ex           (core_i.controller_i.controller_fsm_i.branch_in_ex),

      .mie_q                  (core_i.cs_registers_i.mie_q),
      .dcsr_q                 (core_i.cs_registers_i.dcsr_q),
      .depc_q                 (core_i.cs_registers_i.dpc_q),
      .depc_n                 (core_i.cs_registers_i.dpc_n),
      .mcause_q               (core_i.cs_registers_i.mcause_q),
      .mtvec                  (core_i.cs_registers_i.mtvec_q),
      .mepc_q                 (core_i.cs_registers_i.mepc_q),
      .tdata1                 (core_i.cs_registers_i.tdata1_q),
      .tdata2                 (core_i.cs_registers_i.tdata2_q),
      .mcountinhibit_q        (core_i.cs_registers_i.mcountinhibit_q),
      .mcycle                 (core_i.cs_registers_i.mhpmcounter_q[0]),
      .minstret               (core_i.cs_registers_i.mhpmcounter_q[2]),
      .csr_we_int             (core_i.cs_registers_i.csr_we_int),

      // TODO: review this change from CV32E40S_HASH f6196bf to a26b194. It should be logically equivalent.
      //assign debug_cov_assert_if.inst_ret = core_i.cs_registers_i.inst_ret;
      // First attempt: this causes unexpected failures of a_minstret_count
      //assign debug_cov_assert_if.inst_ret = (core_i.id_valid &
      //                                       core_i.is_decoding);
      // Second attempt: (based on OK input).  This passes, but maybe only because p_minstret_count
      //                                       is the only property sensitive to inst_ret. Will
      //                                       this work in the general case?
      .inst_ret               (core_i.ctrl_fsm.mhpmevent.minstret),
      .csr_access             (core_i.ex_wb_pipe.csr_en),
      .csr_op                 (core_i.ex_wb_pipe.csr_op),
      .csr_addr               (core_i.ex_wb_pipe.csr_addr),
      .irq_ack_o              (core_i.irq_ack),
      .irq_id_o               (core_i.irq_id),
      .dm_halt_addr_i         (core_i.dm_halt_addr_i),
      .dm_exception_addr_i    (core_i.dm_exception_addr_i),
      .core_sleep_o           (core_i.core_sleep_o),
      .irq_i                  (core_i.irq_i),
      .pc_set                 (core_i.ctrl_fsm.pc_set),
      .boot_addr_i            (core_i.boot_addr_i),

      .rvfi_valid             (rvfi_i.rvfi_valid),
      .rvfi_insn              (rvfi_i.rvfi_insn),
      .rvfi_intr              (rvfi_i.rvfi_intr),
      .rvfi_dbg               (rvfi_i.rvfi_dbg),
      .rvfi_dbg_mode          (rvfi_i.rvfi_dbg_mode),
      .rvfi_pc_wdata          (rvfi_i.rvfi_pc_wdata),
      .rvfi_pc_rdata          (rvfi_i.rvfi_pc_rdata),
      .rvfi_csr_dpc_rdata     (rvfi_i.rvfi_csr_dpc_rdata),
      .rvfi_csr_mepc_wdata    (rvfi_i.rvfi_csr_mepc_wdata),
      .rvfi_csr_mepc_wmask    (rvfi_i.rvfi_csr_mepc_wmask),
      .rvfi_csr_mepc_rdata    (rvfi_i.rvfi_csr_mepc_rdata),



      .is_wfi                 (),
      .in_wfi                 (),
      .dpc_will_hit           (),
      .addr_match             (),
      .is_ebreak              (),
      .is_cebreak             (),
      .is_dret                (),
      .is_mulhsu              (),
      .pending_enabled_irq    (),

      .*
    );


    bind cv32e40s_wrapper
      uvmt_cv32e40s_support_logic_if support_logic_if ();

    // TODO find a better way
    assign dut_wrap.cv32e40s_wrapper_i.support_logic_if.ctrl_fsm_o_i   = dut_wrap.cv32e40s_wrapper_i.core_i.controller_i.controller_fsm_i.ctrl_fsm_o;
    assign dut_wrap.cv32e40s_wrapper_i.support_logic_if.data_bus_req_i = dut_wrap.cv32e40s_wrapper_i.core_i.m_c_obi_data_if.s_req.req;
    assign dut_wrap.cv32e40s_wrapper_i.support_logic_if.data_bus_gnt_i = dut_wrap.cv32e40s_wrapper_i.core_i.m_c_obi_data_if.s_gnt.gnt;
    assign dut_wrap.cv32e40s_wrapper_i.support_logic_if.clk_i          = dut_wrap.cv32e40s_wrapper_i.core_i.clk_i;
    assign dut_wrap.cv32e40s_wrapper_i.support_logic_if.rst_ni         = dut_wrap.cv32e40s_wrapper_i.core_i.rst_ni;


    bind cv32e40s_pmp :
      uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.if_stage_i.mpu_i.pmp.pmp_i
      uvmt_cv32e40s_pmp_assert#(
        .PMP_GRANULARITY(PMP_GRANULARITY),
        .PMP_NUM_REGIONS(PMP_NUM_REGIONS),
        .IS_INSTR_SIDE(1'b1),
        .MSECCFG_RESET_VAL(cv32e40s_pkg::MSECCFG_DEFAULT)
      )
      u_pmp_assert_if_stage(.rst_n (clknrst_if.reset_n),
                            .obi_req (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_req_o),
                            .obi_addr (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_addr_o),
                            .obi_gnt (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.instr_gnt_i),
                            .rvfi_valid (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_valid),
                            .rvfi_pc_rdata (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_pc_rdata),
                            .*);

    bind  cv32e40s_pmp :
      uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.load_store_unit_i.mpu_i.pmp.pmp_i
      uvmt_cv32e40s_pmp_assert#(
        .PMP_GRANULARITY(PMP_GRANULARITY),
        .PMP_NUM_REGIONS(PMP_NUM_REGIONS),
        .IS_INSTR_SIDE(1'b0),
        .MSECCFG_RESET_VAL(cv32e40s_pkg::MSECCFG_DEFAULT)
      )
      u_pmp_assert_lsu(.rst_n (clknrst_if.reset_n),
                       .obi_req (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_req_o),
                       .obi_addr (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_addr_o),
                       .obi_gnt (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.core_i.data_gnt_i),
                       .rvfi_valid (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_valid),
                       .rvfi_pc_rdata (uvmt_cv32e40s_tb.dut_wrap.cv32e40s_wrapper_i.rvfi_i.rvfi_pc_rdata),
                       .*);

    bind  dut_wrap.cv32e40s_wrapper_i.rvfi_i
      uvmt_cv32e40s_pmprvfi_assert #(
        .PMP_GRANULARITY (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_GRANULARITY),
        .PMP_NUM_REGIONS (uvmt_cv32e40s_pkg::CORE_PARAM_PMP_NUM_REGIONS)
      ) pmprvfi_assert_i (
        .rvfi_mem_addr  (rvfi_mem_addr [31:0]),
        .rvfi_mem_wmask (rvfi_mem_wmask[ 3:0]),
        .rvfi_mem_rmask (rvfi_mem_rmask[ 3:0]),
        .*
      );

    bind cv32e40s_wrapper uvmt_cv32e40s_support_logic u_support_logic(.rvfi(rvfi_instr_if_0_i),
                                                                      .support_if(support_logic_if)
                                                                      );

    bind cv32e40s_wrapper uvmt_cv32e40s_debug_assert u_debug_assert(.cov_assert_if(debug_cov_assert_if));

    bind cv32e40s_wrapper uvmt_cv32e40s_zc_assert u_zc_assert(.rvfi(rvfi_instr_if_0_i),
                                                              .support_if(support_logic_if)
                                                              );


    //uvmt_cv32e40s_rvvi_handcar u_rvvi_handcar();
    /**
    * ISS WRAPPER instance:
    */
    `ifndef FORMAL
      uvmt_cv32e40s_iss_wrap  #(
                                .ID (0),
                                .ROM_START_ADDR('h0),
                                .ROM_BYTE_SIZE('h0),
                                .RAM_BYTE_SIZE('h1_0000_0000)
                               )
                               iss_wrap ( .clk_period(clknrst_if.clk_period),
                                          .clknrst_if(clknrst_if_iss)
                                 );

      assign clknrst_if_iss.reset_n = clknrst_if.reset_n;
    `endif

   /**
    * Test bench entry point.
    */
   `ifndef FORMAL // Formal ignores initial blocks, avoids unnecessary warning
   initial begin : test_bench_entry_point

     // Specify time format for simulation (units_number, precision_number, suffix_string, minimum_field_width)
     $timeformat(-9, 3, " ns", 8);

     // Add interfaces handles to uvm_config_db
     uvm_config_db#(virtual uvma_isacov_if              )::set(.cntxt(null), .inst_name("*.env.isacov_agent"),           .field_name("vif"),           .value(isacov_if));
     uvm_config_db#(virtual uvma_debug_if               )::set(.cntxt(null), .inst_name("*.env.debug_agent"),            .field_name("vif"),           .value(debug_if));
     uvm_config_db#(virtual uvma_clknrst_if             )::set(.cntxt(null), .inst_name("*.env.clknrst_agent"),          .field_name("vif"),           .value(clknrst_if));
     uvm_config_db#(virtual uvma_interrupt_if           )::set(.cntxt(null), .inst_name("*.env.interrupt_agent"),        .field_name("vif"),           .value(interrupt_if));
     uvm_config_db#(virtual uvma_clic_if                )::set(.cntxt(null), .inst_name("*.env.clic_agent"),             .field_name("vif"),           .value(clic_if));
     uvm_config_db#(virtual uvma_obi_memory_if          )::set(.cntxt(null), .inst_name("*.env.obi_memory_instr_agent"), .field_name("vif"),           .value(obi_instr_if_i) );
     uvm_config_db#(virtual uvma_obi_memory_if          )::set(.cntxt(null), .inst_name("*.env.obi_memory_data_agent"),  .field_name("vif"),           .value(obi_data_if_i) );
     uvm_config_db#(virtual uvma_fencei_if              )::set(.cntxt(null), .inst_name("*.env.fencei"),                 .field_name("vif"),           .value(fencei_if_i));
     uvm_config_db#(virtual uvma_rvfi_instr_if          )::set(.cntxt(null), .inst_name("*.env.rvfi_agent"),             .field_name("instr_vif0"),    .value(dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i));
     uvm_config_db#(virtual uvma_fencei_if              )::set(.cntxt(null), .inst_name("*.env.fencei_agent"),           .field_name("fencei_vif"),    .value(fencei_if_i)  );
     uvm_config_db#(virtual uvmt_cv32e40s_vp_status_if  )::set(.cntxt(null), .inst_name("*"),                            .field_name("vp_status_vif"), .value(vp_status_if) );
     uvm_config_db#(virtual uvma_interrupt_if           )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("intr_vif"),      .value(interrupt_if) );
     uvm_config_db#(virtual uvma_clic_if                )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("clic_vif"),      .value(clic_if) );
     uvm_config_db#(virtual uvma_debug_if               )::set(.cntxt(null), .inst_name("*.env"),                        .field_name("debug_vif"),     .value(debug_if)     );
//     uvm_config_db#(virtual uvmt_cv32e40s_debug_cov_assert_if)::set(.cntxt(null), .inst_name("*.env"),                 .field_name("debug_cov_vif"),    .value(debug_cov_assert_if));
     `RVFI_CSR_UVM_CONFIG_DB_SET(marchid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcountinhibit)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstatus)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mstatush)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcounteren)
     `RVFI_CSR_UVM_CONFIG_DB_SET(menvcfg)
     `RVFI_CSR_UVM_CONFIG_DB_SET(menvcfgh)
     `RVFI_CSR_UVM_CONFIG_DB_SET(misa)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mtvec)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mtval)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mvendorid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mscratch)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mepc)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcause)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mip)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mie)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhartid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mimpid)
     `RVFI_CSR_UVM_CONFIG_DB_SET(minstret)
     `RVFI_CSR_UVM_CONFIG_DB_SET(minstreth)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcycle)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mcycleh)

     `RVFI_CSR_UVM_CONFIG_DB_SET(dcsr)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dpc)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dscratch0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(dscratch1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tselect)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tdata3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(tinfo)

     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpcfg15)

     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr0)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr1)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr2)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr31)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr32)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr33)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr34)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr35)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr36)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr37)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr38)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr39)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr40)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr41)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr42)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr43)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr44)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr45)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr46)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr47)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr48)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr49)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr50)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr51)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr52)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr53)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr54)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr55)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr56)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr57)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr58)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr59)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr60)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr61)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr62)
     `RVFI_CSR_UVM_CONFIG_DB_SET(pmpaddr63)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmevent31)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter3)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter4)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter5)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter6)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter7)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter8)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter9)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter10)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter11)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter12)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter13)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter14)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter15)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter16)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter17)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter18)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter19)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter20)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter21)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter22)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter23)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter24)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter25)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter26)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter27)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter28)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter29)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter30)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter31)

     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter3h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter4h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter5h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter6h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter7h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter8h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter9h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter10h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter11h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter12h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter13h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter14h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter15h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter16h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter17h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter18h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter19h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter20h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter21h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter22h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter23h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter24h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter25h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter26h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter27h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter28h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter29h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter30h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mhpmcounter31h)
     `RVFI_CSR_UVM_CONFIG_DB_SET(mconfigptr)

     uvm_config_db#(virtual RVVI_state#(.ILEN(uvme_cv32e40s_pkg::ILEN),
                                        .XLEN(uvme_cv32e40s_pkg::XLEN)
                                        ))::set(.cntxt(null), .inst_name("*.env.rvvi_agent"), .field_name("state_vif"), .value(iss_wrap.cpu.state));
     uvm_config_db#(virtual RVVI_control                )::set(.cntxt(null), .inst_name("*.env.rvvi_agent"), .field_name("control_vif"), .value(iss_wrap.cpu.control));
     uvm_config_db#(virtual RVVI_bus                    )::set(.cntxt(null), .inst_name("*.env.rvvi_agent"), .field_name("ovpsim_bus_vif"), .value(iss_wrap.bus));
     uvm_config_db#(virtual RVVI_io                     )::set(.cntxt(null), .inst_name("*.env.rvvi_agent"), .field_name("ovpsim_io_vif"), .value(iss_wrap.io));
     uvm_config_db#(virtual RVVI_memory                 )::set(.cntxt(null), .inst_name("*.env.rvvi_agent"), .field_name("ovpsim_mem_vif"), .value(iss_wrap.ram.memory));
     uvm_config_db#(virtual uvmt_cv32e40s_vp_status_if      )::set(.cntxt(null), .inst_name("*"), .field_name("vp_status_vif"),       .value(vp_status_if)      );
     uvm_config_db#(virtual uvme_cv32e40s_core_cntrl_if     )::set(.cntxt(null), .inst_name("*"), .field_name("core_cntrl_vif"),      .value(core_cntrl_if)     );
     uvm_config_db#(virtual uvmt_cv32e40s_core_status_if    )::set(.cntxt(null), .inst_name("*"), .field_name("core_status_vif"),     .value(core_status_if)    );
     uvm_config_db#(virtual uvmt_cv32e40s_debug_cov_assert_if)::set(.cntxt(null), .inst_name("*.env"), .field_name("debug_cov_vif"),.value(dut_wrap.cv32e40s_wrapper_i.debug_cov_assert_if));
     uvm_config_db#(virtual uvmt_cv32e40s_support_logic_if)::set(.cntxt(null), .inst_name("*.env"), .field_name("support_logic_vif"),.value(dut_wrap.cv32e40s_wrapper_i.support_logic_if));

     // Make the DUT Wrapper Virtual Peripheral's status outputs available to the base_test
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("tp"),     .value(1'b0)        );
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("tf"),     .value(1'b0)        );
     uvm_config_db#(bit      )::set(.cntxt(null), .inst_name("*"), .field_name("evalid"), .value(1'b0)        );
     uvm_config_db#(bit[31:0])::set(.cntxt(null), .inst_name("*"), .field_name("evalue"), .value(32'h00000000));

	 // DUT and ENV parameters
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_INSTR_ADDR_WIDTH"),  .value(ENV_PARAM_INSTR_ADDR_WIDTH) );
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_INSTR_DATA_WIDTH"),  .value(ENV_PARAM_INSTR_DATA_WIDTH) );
     uvm_config_db#(int)::set(.cntxt(null), .inst_name("*"), .field_name("ENV_PARAM_RAM_ADDR_WIDTH"),    .value(ENV_PARAM_RAM_ADDR_WIDTH)   );

     // Run test
     uvm_top.enable_print_topology = 0; // ENV coders enable this as a debug aid
     uvm_top.finish_on_completion  = 1;
     uvm_top.run_test();
   end : test_bench_entry_point
   `endif

   assign core_cntrl_if.clk = clknrst_if.clk;
  `ifndef  FORMAL
     assign iss_wrap.cpu.io.nmi_addr = ({dut_wrap.cv32e40s_wrapper_i.rvfi_csr_mtvec_if_0_i.rvfi_csr_rdata[31:2], 2'b00}) + 32'h3c;
  `endif

   // Informational print message on loading of OVPSIM ISS to benchmark some elf image loading times
   // OVPSIM runs its initialization at the #1ns timestamp, and should dominate the initial startup time
   longint start_ovpsim_init_time;
   longint end_ovpsim_init_time;
   `ifndef FORMAL // Formal ignores initial blocks, avoids unnecessary warning
   initial begin
      if (!$test$plusargs("DISABLE_OVPSIM")) begin
        #0.9ns;
        `uvm_info("OVPSIM", $sformatf("Start benchmarking OVPSIM initialization"), UVM_LOW)
        start_ovpsim_init_time = svlib_pkg::sys_dayTime();
        #1.1ns;
        end_ovpsim_init_time = svlib_pkg::sys_dayTime();
        `uvm_info("OVPSIM", $sformatf("Initialization time: %0d seconds", end_ovpsim_init_time - start_ovpsim_init_time), UVM_LOW)
      end
    end
   `endif

   //TODO verify these are correct with regards to isacov function
   `ifndef FORMAL // events ignored for formal - this avoids unnecessary warning
   always @(dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i.rvfi_valid) -> isacov_if.retire;
   `endif
   assign isacov_if.instr = dut_wrap.cv32e40s_wrapper_i.rvfi_instr_if_0_i.rvfi_insn;
   //assign isacov_if.is_compressed = dut_wrap.cv32e40s_wrapper_i.tracer_i.insn_compressed;

   // Capture the test status and exit pulse flags
   // TODO: put this logic in the vp_status_if (makes it easier to pass to ENV)
   always @(posedge clknrst_if.clk) begin
     if (!clknrst_if.reset_n) begin
       tp     <= 1'b0;
       tf     <= 1'b0;
       evalid <= 1'b0;
       evalue <= 32'h00000000;
     end
     else begin
       if (vp_status_if.tests_passed) begin
         tp <= 1'b1;
         uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("tp"), .value(1'b1));
       end
       if (vp_status_if.tests_failed) begin
         tf <= 1'b1;
         uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("tf"), .value(1'b1));
       end
       if (vp_status_if.exit_valid) begin
         evalid <= 1'b1;
         uvm_config_db#(bit)::set(.cntxt(null), .inst_name("*"), .field_name("evalid"), .value(1'b1));
       end
       if (vp_status_if.exit_valid) begin
         evalue <= vp_status_if.exit_value;
         uvm_config_db#(bit[31:0])::set(.cntxt(null), .inst_name("*"), .field_name("evalue"), .value(vp_status_if.exit_value));
       end
     end
   end


   /**
    * End-of-test summary printout.
    */
   `ifndef FORMAL // Formal ignores final blocks, this avoids unnecessary warning
   final begin: end_of_test
      string             summary_string;
      uvm_report_server  rs;
      int                err_count;
      int                warning_count;
      int                fatal_count;
      static bit         sim_finished = 0;

      static string  red   = "\033[31m\033[1m";
      static string  green = "\033[32m\033[1m";
      static string  reset = "\033[0m";

      rs            = uvm_top.get_report_server();
      err_count     = rs.get_severity_count(UVM_ERROR);
      warning_count = rs.get_severity_count(UVM_WARNING);
      fatal_count   = rs.get_severity_count(UVM_FATAL);

      void'(uvm_config_db#(bit)::get(null, "", "sim_finished", sim_finished));

      $display("\n%m: *** Test Summary ***\n");

      if (sim_finished && (err_count == 0) && (fatal_count == 0)) begin
         $display("    PPPPPPP    AAAAAA    SSSSSS    SSSSSS   EEEEEEEE  DDDDDDD     ");
         $display("    PP    PP  AA    AA  SS    SS  SS    SS  EE        DD    DD    ");
         $display("    PP    PP  AA    AA  SS        SS        EE        DD    DD    ");
         $display("    PPPPPPP   AAAAAAAA   SSSSSS    SSSSSS   EEEEE     DD    DD    ");
         $display("    PP        AA    AA        SS        SS  EE        DD    DD    ");
         $display("    PP        AA    AA  SS    SS  SS    SS  EE        DD    DD    ");
         $display("    PP        AA    AA   SSSSSS    SSSSSS   EEEEEEEE  DDDDDDD     ");
         $display("    ----------------------------------------------------------");
         if (warning_count == 0) begin
           $display("                        SIMULATION PASSED                     ");
         end
         else begin
           $display("                 SIMULATION PASSED with WARNINGS              ");
         end
         $display("    ----------------------------------------------------------");
      end
      else begin
         $display("    FFFFFFFF   AAAAAA   IIIIII  LL        EEEEEEEE  DDDDDDD       ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FFFFF     AAAAAAAA    II    LL        EEEEE     DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA    II    LL        EE        DD    DD      ");
         $display("    FF        AA    AA  IIIIII  LLLLLLLL  EEEEEEEE  DDDDDDD       ");

         if (sim_finished == 0) begin
            $display("    --------------------------------------------------------");
            $display("                   SIMULATION FAILED - ABORTED              ");
            $display("    --------------------------------------------------------");
         end
         else begin
            $display("    --------------------------------------------------------");
            $display("                       SIMULATION FAILED                    ");
            $display("    --------------------------------------------------------");
         end
      end
   end
   `endif

endmodule : uvmt_cv32e40s_tb
`default_nettype wire

`endif // __UVMT_CV32E40S_TB_SV__
