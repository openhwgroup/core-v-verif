// Copyright 2023 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// -------------------------------------------------------------------
// This file holds constants related to the ISA
// -------------------------------------------------------------------

`ifndef __ISA_CONSTANTS__
`define __ISA_CONSTANTS__

parameter CLIC_ID_WIDTH = 5;
parameter DEFAULT_XLEN = 32;

`endif // __ISA_CONSTANTS__
