// Copyright 2020 OpenHW Group
// Copyright 2020 Datum Technology Corporation
// Copyright 2024 Dolphin Design
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//

// This file specifies all interfaces used by the CV32E40P test bench (uvmt_cv32e40p_tb), related to DUT control.
// Most interfaces support tasks to allow control by the ENV or test cases.

`ifndef __UVMT_CV32E40P_TB_DUT_IFS_SV__
`define __UVMT_CV32E40P_TB_DUT_IFS_SV__



/**
 * clocks and reset
 */
 interface uvmt_cv32e40p_clk_gen_if (output logic core_clock, output logic core_reset_n);

    import uvm_pkg::*;

    bit       start_clk               = 0;
    // TODO: get the uvme_cv32e40p_* values from random ENV CFG members.
    realtime  core_clock_period       = 1500ps; // uvme_cv32e40p_clk_period * 1ps;
    realtime  reset_deassert_duration = 7400ps; // uvme_cv32e40p_reset_deassert_duarion * 1ps;
    realtime  reset_assert_duration   = 7400ps; // uvme_cv32e40p_reset_assert_duarion * 1ps;


    /**
     * Generates clock and reset signals.
     * If reset_n comes up de-asserted (1'b1), wait a bit, then assert, then de-assert
     * Otherwise, leave reset asserted, wait a bit, then de-assert.
     */
    initial begin
       core_clock   = 0; // uvme_cv32e40p_clk_initial_value;
       core_reset_n = 0; // uvme_cv32e40p_reset_initial_value;
       wait (start_clk);
       fork
          forever begin
             #(core_clock_period/2) core_clock = ~core_clock;
          end
          begin
            if (core_reset_n == 1'b1) #(reset_deassert_duration);
            core_reset_n = 1'b0;
            #(reset_assert_duration);
            core_reset_n = 1'b1;
          end
       join_none
    end

    /**
     * Sets clock period in ps.
     */
    function static void set_clk_period ( real clk_period );
       core_clock_period = clk_period * 1ps;
    endfunction : set_clk_period

    /** Triggers the generation of clk. */
    function static void start();
       start_clk = 1;
       `uvm_info("CLK_GEN_IF", "uvmt_cv32e40p_clk_gen_if.start() called", UVM_NONE)
    endfunction : start

 endinterface : uvmt_cv32e40p_clk_gen_if

 /**
  * Status information generated by the Virtual Peripherals in the DUT WRAPPER memory.
  */
 interface uvmt_cv32e40p_vp_status_if (
                                   output reg        tests_passed,
                                   output reg        tests_failed,
                                   output reg        exit_valid,
                                   output reg [31:0] exit_value
                                  );

   import uvm_pkg::*;

   // TODO: X/Z checks
   initial begin
   end

 endinterface : uvmt_cv32e40p_vp_status_if



 /**
  * Core status signals.
  */
 interface uvmt_cv32e40p_core_status_if (
                                     input  wire        core_busy,
                                     input  logic       sec_lvl
                                    );

   import uvm_pkg::*;

 endinterface : uvmt_cv32e40p_core_status_if


 // Interface to debug assertions and covergroups
interface uvmt_cv32e40p_debug_cov_assert_if
   import cv32e40p_pkg::*;
   (
   input  clk_i,
   input  rst_ni,

   // Core inputs
   input         fetch_enable_i, // external core fetch enable

   // External interrupt interface
   input  [31:0] irq_i,
   input         irq_ack_o,
   input  [4:0]  irq_id_o,
   input  [31:0] mie_q,

   // Instruction fetch stage
   input         if_stage_instr_rvalid_i, // Instruction word is valid
   input  [31:0] if_stage_instr_rdata_i, // Instruction word data

   // Instruction ID stage (determines executed instructions)
   input         id_stage_instr_valid_i, // instruction word is valid
   input  [31:0] id_stage_instr_rdata_i, // Instruction word data
   input         id_stage_is_compressed,
   input  [31:0] id_stage_pc, // Program counter in decode
   input  [31:0] if_stage_pc, // Program counter in fetch
   input         is_decoding,
   input         branch_taken_ex_i,
   input         data_err_i,
   input         is_fetch_failed_i,
   input         id_valid,
   input wire ctrl_state_e  ctrl_fsm_cs,            // Controller FSM states with debug_req
   input         illegal_insn_i,
   input         illegal_insn_q, // output from controller
   input         ecall_insn_i,

   input  [31:0] boot_addr_i,

   input         rvfi_valid,
   input  [31:0] rvfi_insn,
   input         apu_req,
   input         apu_gnt,
   input         apu_busy,

   // Debug signals
   input         debug_req_i, // From controller
   input         debug_mode_q, // From controller
   input  [31:0] dcsr_q, // From controller
   input  [31:0] depc_q, // From cs regs
   input  [31:0] depc_n, //
   input  [31:0] dm_halt_addr_i,
   input  [31:0] dm_exception_addr_i,

   input  [5:0]  mcause_q,
   input  [31:0] mtvec,
   input  [31:0] mepc_q,
   input  [31:0] tdata1,
   input  [31:0] tdata2,
   input  trigger_match_i,

   // Counter related input from cs_registers
   input  [31:0] mcountinhibit_q,
   input  [63:0] mcycle,
   input  [63:0] minstret,
   input  inst_ret,
   // WFI Interface
   input  core_sleep_o,

   input  fence_i,

   input  csr_access,
   input  [1:0] csr_op,
   input  [1:0] csr_op_dec,
   input  [11:0] csr_addr,
   input  csr_we_int,

   output logic is_wfi,
   output logic in_wfi,
   output logic dpc_will_hit,
   output logic addr_match,
   output logic is_ebreak,
   output logic is_cebreak,
   output logic is_dret,
   output logic is_mulhsu,
   output logic [31:0] pending_enabled_irq,
   input  pc_set,
   input  branch_in_decode
);

 clocking mon_cb @(posedge clk_i);
   input #1step
   fetch_enable_i,

   irq_i,
   irq_ack_o,
   irq_id_o,
   mie_q,

   if_stage_instr_rvalid_i,
   if_stage_instr_rdata_i,

   id_stage_instr_valid_i,
   id_stage_instr_rdata_i,
   id_stage_is_compressed,
   id_stage_pc,
   if_stage_pc,
   is_decoding,
   branch_taken_ex_i,
   is_fetch_failed_i,
   id_valid,
   ctrl_fsm_cs,
   illegal_insn_i,
   illegal_insn_q,
   ecall_insn_i,
   boot_addr_i,
   rvfi_valid,
   rvfi_insn,
   apu_req,
   apu_gnt,
   apu_busy,
   debug_req_i,
   debug_mode_q,
   dcsr_q,
   depc_q,
   depc_n,
   dm_halt_addr_i,
   dm_exception_addr_i,
   mcause_q,
   mtvec,
   mepc_q,
   tdata1,
   tdata2,
   trigger_match_i,
   fence_i,
   mcountinhibit_q,
   mcycle,
   minstret,
   inst_ret,

   core_sleep_o,
   csr_access,
   csr_op,
   csr_op_dec,
   csr_addr,
   is_wfi,
   in_wfi,
   dpc_will_hit,
   addr_match,
   is_ebreak,
   is_cebreak,
   is_dret,
   is_mulhsu,
   pending_enabled_irq,
   pc_set,
   branch_in_decode;
 endclocking : mon_cb

endinterface : uvmt_cv32e40p_debug_cov_assert_if




`endif // __UVMT_CV32E40P_TB_DUT_IFS_SV__
