// Copyright 2024 OpenHW Group
// SPDX-License-Identifier: Apache-2.0 WITH SHL-210
`ifndef __UVMA_CV32E40P_COV_MODEL_MACROS_SV__
`define __UVMA_CV32E40P_COV_MODEL_MACROS_SV__

// Place any CV32E40P coverage model specific macros here...

`endif // __UVMA_CV32E40P_COV_MODEL_MACROS_SV__