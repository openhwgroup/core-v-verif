// ----------------------------------------------------------------
// ----------------------------------------------------------------------------
//                                CEA - LETI
//    Reproduction and Communication of this document is strictly prohibited
//      unless specifically authorized in writing by CEA - LETI.
// ----------------------------------------------------------------------------
//                        LETI / DACLE / LISAN
// ----------------------------------------------------------------------------
//
//
//  File        :
//  Entity      :
//
//  Description :
//
//
//  Copyright (C) 2019 CEA-Leti
//  Author      : $authorname : PERBOST Nicolas $ $authoremail : nicolas.perbost.fr $
//
//  Id          : $Id: ebc1c90d292c16718a5f425063aa10baa9553215 $
//  Date        : $Date : Tue Mar 5 17:22:29 2019 +0100 $
//
// ----------------------------------------------------------------------------

package test_pkg;

    import uvm_pkg::*;
    import uvma_axi_pkg::*;
    import dut_env_pkg::*;
    `include "uvm_macros.svh";
    `include "base_test_c.svh";
    `include "bursty_test_c.svh";


endpackage : test_pkg


