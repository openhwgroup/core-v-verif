// Add your custom extensions, you can list all your local extended SV files here
`include "isa/custom/cv32e40p_defines.svh"
