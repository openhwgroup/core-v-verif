//
// Copyright 2023 OpenHW Group
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//

`ifndef __UVMT_CV32E40S_BASE_TEST_CONSTRAINT_WORKAROUNDS_SV__
`define __UVMT_CV32E40S_BASE_TEST_CONSTRAINT_WORKAROUNDS_SV__


// This file should be empty by the end of the project

`endif // __UVMT_CV32E40S_BASE_TEST_CONSTRAINT_WORKAROUNDS_SV__
