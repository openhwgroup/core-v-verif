// Copyright 2023 Silicon Labs, Inc.
//
// Licensed under the Solderpad Hardware Licence, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     https://solderpad.org/licenses/
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0

`ifndef __ISA_DECODER_PKG__
`define __ISA_DECODER_PKG__


package isa_decoder_pkg;
  `include "isa_constants.sv"
  `include "isa_typedefs_csr.sv"
  `include "isa_typedefs.sv"
  `include "isa_decoder.sv"
endpackage

`endif // __ISA_DECODER_PKG__

