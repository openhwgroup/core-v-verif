/*
 * Copyright 2023 Dolphin Design
 * SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 */

`DEFINE_FP_IN_X_INSTR(FMADD_S,   R4_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FMSUB_S,   R4_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FNMSUB_S,  R4_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FNMADD_S,  R4_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FADD_S,    R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FSUB_S,    R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FMUL_S,    R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FDIV_S,    R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FSQRT_S,   I_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FSGNJ_S,   R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FSGNJN_S,  R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FSGNJX_S,  R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FMIN_S,    R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FMAX_S,    R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FCVT_W_S,  I_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FCVT_WU_S, I_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FEQ_S,     R_FORMAT, COMPARE, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FLT_S,     R_FORMAT, COMPARE, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FLE_S,     R_FORMAT, COMPARE, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FCLASS_S,  R_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FCVT_S_W,  I_FORMAT, ARITHMETIC, RV32ZFINX)
`DEFINE_FP_IN_X_INSTR(FCVT_S_WU, I_FORMAT, ARITHMETIC, RV32ZFINX)
